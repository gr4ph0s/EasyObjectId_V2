MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$       "	�fhc�fhc�fhc�k:��ehc��Ȥ�ghc�k:��ehc�k:��mhc�k:��bhc껗��dhc�fhb�@hc�C��@hc�C��ghc�k:��ghc�C��ghc�Richfhc�                PE  L ���Y        � !    B      e                                 �         @                   pA L   �A <    ` �                   p �  �  8                           �: @              �                           .text   I                        `.rdata  �$      &                @  @.data   �   P     :             @  �.rsrc   �   `     <             @  @.reloc  �   p     >             @  B                                                                                                                                                                                                                                                                                                                                h �  Y������ ����U�h�v  Y����̡ UV�r�2�@����� VQ���   �Ѓ�^��������������U�� UV��V�@�@�С Uj j��u�@V�@�Ѓ���^]� �������������� �������������� �������������U���EV����5t
V�l ����^]� ������������̡ UVW���    �w@�G   �G    �G    �G    �G    �G    �G    �G     �G$    �G(    �G,    �G4   �G8   �G<    �@V�@�С Uj j�h4�@V�@�Ѓ��GP_   �GT  4B���GX    �G\    �G`   �Gd   �Gh    _^����U��SV��W�}�s@V�o��oG�C�oG �C �G0�C0�G4�C4�G8�C8�G<�C<� U�@�@�С UV�H�G@P�A�ЋGP���CP�GT�CT�GX�CX�G\�C\�G`�C`�Gd�Cd�Gh_�Ch��^[]� ��������U�� UVW��Wh�� ��9�@0� �Ћu�O���G�G    �L6V�   �F8���   ���   �F<���   �F@���   �FD���   �FHP�����ǇH      ��ǇL      _^]� ���U��V����   �Et
V�l ����^]� ��������������U�� USV�ً@WS�@�С US�@$�@D�С U�}SW�@$�@L�С U�sV�@�@�С UV�@$�@D�С UV�H$�GP�AL�ЋG8�KH�C8�� �G<�C<�G@�C@�GD�CD�GHP����_^��[]� ��������̡ US��V�PW��  P�B�С U�{�H���   P�A�С U�wV�@$�@H�С UV�@�@�С UW�@$�@H�С UW�@�@�ЋK����9��t� UQ�@0�@�Ѓ�_^�C    [����������U��V����4�N��t� UQ�@� �Ѓ��F    �E�F    �F    ��5t
V�l ����^]� �����������U��V��N��5��  �E��5t
V�l ����^]� ���������������U��V��N�5�  �E��5t
V�l ����^]� ���������������U��Q�EV��M�F��5�F    �F    �F    �F    �F   ��F�A�ΉF��  �ΉF��  �F ��t���-�  ��^Y]� �����U��V����5�N��t� UQ�@� �Ѓ��F    �E�F    �F    ��5t
V�l ����^]� �����������U��Q�EV��M�F�d5�F    �F    �F    �F    �F   ��F�A�ΉF�u�  �F��t���w�  ��^Y]� ���������������U��V���d5�N��t� UQ�@� �Ѓ��F    �E�F    �F    ��5t
V�l ����^]� �����������U��EVW���G�O�45�G    �G    �G    ��������I�  �u�O�G�{   ��_^]� ���U�� UV���45�P�FXP�B�ЋN����t� UQ�@� �Ѓ��F    �E�F    �F    ��5t
V�l ����^]� �������U��V�uW���o��oF�G�oF �G �F0�G0�F4�G4�F8�G8�F<�G<� U�H�G@P�F@P�A�ЋFP���GP�FT�GT�FX�GX�F\�G\�F`�G`�Fd�Gd�Fh�Gh��_^]� ��������U��V���U  �Et
V�l ����^]� ��������������W���? t=V�wNx,S����� U��Q�@�@�Ѓ���Ny�[^�G    _�^�G    _��G    _���V��> tFW�~Ox"S����� U��Q�@�@�Ѓ���Oy�[�_��t� UQ�@� �Ѓ��    �F    �F    ^��̡ UV��V�@�@�Ѓ���^���������SV��F��X���N;�~yAW�I�+����ρ�  �yI���Au��u	�   +��� Uh�8h�   �H��    P�6��  �ЋЃ���t�N�~_�^���^[� �F_�F��^[� �^^[� ���������U��QV��F�V�H���M�;���   BS�R�+����ˁ�  �yI���Au��u	�   +�ء UWh�8h�   �H����P���  �Ћ�����tM���t)�v���\   �����t� UQ�@� �Ѓ��    �F���>��E��F��_�^[^��]� �F�F��_[^��]� �N^��]� ����U��S�]VW���;�vR����   ��$    ��t � UV�@�@�С UVW�@�@�Ѓ�� UW�@�@�Ѓ�����Ku�_^[]Ë�������~<����t � UV�@�@�С UVW�@�@�Ѓ�� UW�@�@�Ѓ�Ku�_^[]����������������U��V��W���t� UQ�@� �Ѓ��    �}�F    �F    h�8�G�Fh  ��    � UQ�@���  �Ѓ���tH��O�N��Q�7P�� ����u-��F��t� UQ�@� �Ѓ��    �F    �F    �N3�;O_��^]� ����U���EV����9t
V�l ����^]� ��`��` ��`��`��`��`��`��`�����U�� U�@�E    ���   ]�������U��V��N��9��t� UQ�@0�@�Ѓ��E�F    t
V�l ����^]� ��������������U��V��~ �:u� U�v�@4� �Ѓ��E�F    �F    t
V�l ����^]� �������U�� UV���v�H:�@l�@�Ѓ��Et
V�l ����^]� ����������3���������������U��V��~ ��:u� U�v�@P�@�Ѓ��Et
V�l ����^]� �%t �%l U���EV��t%Wh�# �~��7jV�  �EtW�����Y��_��t  �EtV����Y��^]� Vh�   �0 Y��V� ��U��U��u3�@^Ã& �*  h�% �C  �$�% �7  Y3�^�U��QQ�} SVW�)  ��Q���  H��U��Q3�d�   �}��P�;�t3�������u���E�   �=�Utj�  Y�  �5�U� ���u����   �5�U� �؉u�]��;�r\9;t�W� 9t��3� W��� ����5�U�5 ���5�U�E��֋M�9Mu�u9Et���M�u�؉E띃��tV�D YW� ��U��U��U�=�U9}���   3���   3��   �}��   d�   3�����U�P�;�t3�������u��3�F9=�Uj_t	j�  �5h� h� ��U   �  YY��u�h� h� �  Y�=�UY��u3���=�U th�U�  Y��t�uW�u��U��Q3�@_^[��]� U��}u�n  �u�u�u�   ��]� jhh@�L  3�@���u�3ۉ]��}�= P�E���u9=�Q��   ;�t��u8�� ��t�uW�u�Ћ��u����   �uW�u�}������u����   �uW�u��  ���u��u.��u*�uS�u��  �uS�u�>����� ��t	�uS�u�Ѕ�t��uK�uW�u�������#��u�t4�� ��t+�uW�u�Ћ���M�� �E�QP��  YYËe�3ۋ�u�]��E������   ���y  Ëu�� P����Ã=�U t3��Vjj �p YY��V� ��U��U��ujX^Ã& 3�^�jh�@��  �e� �5�U�5 �։E���u�u�L Y�ej�,  Y�e� �5�U�։E��5�U�։E��E�P�E�P�u�5 ��P�  �����}��u��֣�U�u��֣�U�E������   ���  Ë}�j��  Y�U���u�L�����Y���H]�jh�@�  �e� �]�Ë}�ǋu��u�e� O�}x+�u���U��3�@�E��E������   �   � �}�]�u�E��u�uWSV�   �jh�@�  �e� �Mx:�M+M�M�U��E�E�E� �E��E��8csm�t�E�    �E����  �e��E������  � �%$ �%( �%, ������������U��E3�SVW�H<��A�Y�����t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h�@h9& d�    P��SVW�P1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�U����e� �e� �PVW�N�@��  ��;�t��t	�УP�f�E�P�  �E�3E�E�� 1E�� 1E��E�P� �M��E�3M�3M�3�;�u�O�@����u��G  ��ȉP�щP_^��]�VW�X@�X@����t�Ѓ�;�r�_^�VW�`@�`@����t�Ѓ�;�r�_^���%4 �%8 h�Q�   Y�����������h9& d�5    �D$�l$�l$+�SVW�P1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�U���u�u�u�uhz& hP�3   ��]��%< �%@ �%H �%P �%T ;Pu���D   ��%X U��� j�U�#  �u�!  �=U YYuj�	  Yh	 ��
  Y]�U���$  j��   ��tjY�)� S��R��R��R�5�R�=�Rf�Sf�Sf��Rf��Rf�%�Rf�-�R��S�E �S�E�S�E�S�������PR  �S�R� R	 ��R   �R   jXk� ǀR   jXk� �P�L�jX�� �P�L�h� �������]��%\ �%` �%d �% U���It3���]�VQ�M���  P豿  � U���E�P�I$�IH�ы U�A�M�Q�@�Ѓ�3�����^��]������������������������������
  ���������̸   @� ���������+  �   � ���U����VW�}��W�  ��t|���   ��tr��P�F=d� t3Ht&-�� t-&  u*W���  � =�� t=�� uW����  �W���3   � Uj �@��D  �Ћ��   ����t�j�P_�   ^��]� U���t� UVW�u�@L���E�    �E�    �E�    �@�Ћ��   �}����W�vP�R$�}� uZ� U�M�Q�@�@�С U�MЃ��@j j�h44�@Q�С U�M�j0Q�@�@@�С U�M�Q�@�@�Ѓ���  ���   ��P���   �U�R��P� U�M�Q�@�@�С U�M����@j j�hH4�@Q�С U�H�E��RP�E�P���   �Ћ U�����E��IP�I�ы U���A�M�QV�@�С U�M�Q�@�@�С U�M����@Q�@�С U�M����@j j�h\4�@Q�С U�M�Q�@�@�С U���@�M�Q�M�Q�@�С U�MЃ��@�@<�Ћ Uj�j��Q�M�QP�MЋBL�С U�M�Q�@�@�С U�M����@Q�M�Q�@�С U�M����@�@<�Ћ Uj�j��Q�M�QP�M��BL�С U�M�j0Q�@�@@�С U�M�Q�@�@�С U�MЃ��@Q�@�С U�M����@Q�@�С U�M����@Q�@�С U�M����@Q�@�Ѓ��M������M������_^��]� ���������������U���t� UVW�u�@L���E�    �E�    �E�    �@�Ћ��   �}����W�vP�R(�}� uZ� U�M�Q�@�@�С U�MЃ��@j j�h44�@Q�С U�M�j0Q�@�@@�С U�M�Q�@�@�Ѓ���  ���   ��P���   �U�R��P � U�M�Q�@�@�С U�M����@j j�hH4�@Q�С U�H�E��RP�E�P���   �Ћ U�����E��IP�I�ы U���A�M�QV�@�С U�M�Q�@�@�С U�M����@Q�@�С U�M����@j j�h\4�@Q�С U�M�Q�@�@�С U���@�M�Q�M�Q�@�С U�MЃ��@�@<�Ћ Uj�j��Q�M�QP�MЋBL�С U�M�Q�@�@�С U�M����@Q�M�Q�@�С U�M����@�@<�Ћ Uj�j��Q�M�QP�M��BL�С U�M�j0Q�@�@@�С U�M�Q�@�@�С U�MЃ��@Q�@�С U�M����@Q�@�С U�M����@Q�@�С U�M����@Q�@�Ѓ��M��E�    ��t� UQ�@� �Ѓ�_^��]� �V��W�~���R  �~ u!hP  �h ����t
W�������3��F� U�Nj j �@0j j j ���   j j j j4�q�Ѓ�(��u�N�����  _^���������������U���   S�]�E�    VW����u3�_^[��]� �O�  ��t� US�@L�@,�Ѓ��E�    �M��E�    ��h�  ���  � Uj ���   �M�QP�΋B�ЍM��]�  � U�M�Q���   �@8�Ѓ�=d� �3  ��   =n� t�)  ���  ���  =�� ��  j$�G�G*� �h ������t*�WP�E�U�ˋWTP�U��J�  P���������   �!  3����   �  =�� ��  j �G�G� �h ������t͋OH�E�M�OL�M���P��  P���������   ��  j�Gd� �G�� �h ��������  � US�IL�I,�у��F��5���F    �F    �F    �Q  �F�\  =G� ��   ��   =�� ��   =�� ��   h�   �G�G�� �h ������t.�OX�E�   Q��p����m�����p�����P��  P���w����3��E����   ��   � U�M�Q�@�@�Ѓ���   j�G�� �G�� �h ��������   ��谾  �F���5�F    �F    �F    �y  �F�j=%��t�G    �G    �Yj�G   �G  �h ������t2� US�IL�I,�щF����4�F    �F    �F    �3����   � U�E�3�9_P���   �Ë	�у���_^[��]� ������������S��VW�K�$6��t�j�� U�{�H���   P�A�С U�wV�@$�@H�С UV�@�@�С UW�@$�@H�С UW�@�@�Ѓ���9_^[����������U����� U��$�@Vhh4h�   ���   h�   �Ћ�����t�N�$6�0  �3�� U�L$Q�@�@�С U�L$���@j j�h�4�@Q�С U�L$Q�@�@�С U�L$���@j j�h�4�@Q�Ѓ��D$�T$VP���w�  � U���D$P�I�I�ы U���A�L$Q�@�Ѓ���^��]���U��} V��u��  ��u^]� � U�@���   �ЉE���#  � Ujj�Q�NQ��h� ��Ѕ���  � U�v@�M�@�@,�ЋM��� U�@��  �vD�@,�ЋM��� U�@��  �v8�@,�ЋM��� U�@��  �v<�@,�ЋM��� U�@��  �vL�@,�ЋM��� U�@�h  �vP�@,�ЋM��� U�@�M  �vT�@,�ЋM��� U�@�2  �vX�@,�ЋM��� U�@�  �v\�@,�ЋM��� U�@��   �v`�@,�ЋM��� U�@��   �vd�@,�ЋM��� U�@��   �vh�@,�ЋM��� U�@��   �vl�@,�ЋM��� U�@��   �vp�@,�ЋM��� U�@ty�vt�@,�ЋM��� U�@tb�vx�@,�ЋM��� U�@tK�v|�@,�ЋM��� U�@t4���   �@�ЋM��� U�@t���   �@,�ЋM��� Uu)�@�@��3�� U�EP�I���   �у���^]� �P���   P�BL�ЋM��� U�@t����   �@�Ѕ�� U�@u�M����   �@$Q�M�$�ЋM��� U�@�w������   �@�ЋM��� U�@�Y������   �@�ЋM��� U�@�;������   �@�ЋM��� U�@�������   �@�ЋM��� U�@��������   �@�ЋM��� U�@�@������С U�MQ�@���   �Ѓ��E    �   �����U��UV�u���F8�NH�B�U�F<��F@�B�FD�����j ���*���^]� ����̡ UV��j�@V�@�Ѓ���u�����  ��u3�^á Uj �H�FP�A�Ѓ���uj���������tո   ^����������U�� U���   �@V��M�Q�@�С U�M�Q�@$�@D�С U�M�hp6Q�@$�@d�С U�M�Q�@�@�С U�M�Q�@$�@D�С U�M�h�6Q�@$�@d�Ѝ�t������  � U�M�Q�@�@�С U�M�Q�@$�@D�С U�M�Q��t���Q�@$�@L�С U�M�Q�M�Q�@$�@@�С U�M�Q�@�@�С U�M�Q�@$�@D�С U�Mȃ�@�@$Q�M�Q�@L�С U�M�Q�M�Q�@$�@@�С U�M�VQ�@$�@L�С U�M�Q�@$�@H�С U�M�Q�@�@�С U�M�Q�@$�@H�С U�M�Q�@�@�С U��t���Q�@$�@H�С U��t���Q�@�@�С U�M�Q�@$�@H�С U�M�Q�@�@�С U�M�Q�@$�@H�С U�@�M�Q�@�С U��t�����@�@Q�@�С U��t���Q�@$�@D�С U��t���h�6Q�@$�@d�С U��X���Q�@�@�С U��X���Q�@$�@D�С U��X���hp6Q�@$�@d�С U�M�Q�@�@�С U�M�Q�@$�@D�С U�M�h�6Q�@$�@d�Ѝ�<������  � U�M�Q�@�@�С U�M�Q�@$�@D�С U�M�Q�@$�@L��<���Q�С U�M���@�@$Q�M�Q�@@�С U�M�Q�@�@�С U�M�Q�@$�@D�С U�M�Q�M�Q�@$�@L�С U��X���Q�M�Q�@$�@@�С U�M�Q�@�@�С U�M�Q�@$�@D�С U�M�Q�M�Q�@$�@L�С U��t���Q�M�Q�@$�@@�С U�H$�FP�E�P�AL�С U�M��@�@$�@HQ�С U�M�Q�@�@�С U�M�Q�@$�@H�С U�M�Q�@�@�С U�M�Q�@$�@H�С U�M�Q�@�@�С U��<���Q�@$�@H�С U��<���Q�@�@�С U�M�Q�@$�@H�С U�M�Q�@�@�С U��X���Q�@$�@H�С U��X���Q�@�@�С U��t���Q�@$�@H�С U��t���Q�@�@�Ѓ�8^��]��U����� U�� �@VW��@jV�Ѓ���u����  ��t'� U�~j W�@�@�Ѓ���uj��������u3�_^��]á U�@���   �ЉD$����  � UjjW�Q��h� ��Ѕ���  � U�L$Q�@�@�С U�L$���@Q�L$���   �Ѕ��  �D$�L$�F@� UQ�L$�@���   �Ѕ���  �D$�L$�FD� UQ�L$�@���   �Ѕ���  �D$�L$�F<� UQ�L$�@���   �Ѕ���  �D$�L$�F8� UQ�L$�@���   �Ѕ��y  �D$�L$�FL� UQ�L$�@���   �Ѕ��Q  �D$�L$�FP� UQ�L$�@���   �Ѕ��)  �D$�L$�FT� UQ�L$�@���   �Ѕ��  �D$�L$�FX� UQ�L$�@���   �Ѕ���  �D$�L$�F\� UQ�L$�@���   �Ѕ���  �D$�L$�F`� UQ�L$�@���   �Ѕ���  �D$�L$�Fd� UQ�L$�@���   �Ѕ��a  �D$�L$�Fh� UQ�L$�@���   �Ѕ��9  �D$�L$�Fl� UQ�L$�@���   �Ѕ��  �D$�L$�Fp� UQ�L$�@���   �Ѕ���  �D$�L$�Ft� UQ�L$�@���   �Ѕ���  �D$�L$�Fx� UQ�L$�@���   �Ѕ���  �D$�L$�F|� UQ�L$�@�@p�Ѕ��t  �D$�L$���   � UQ�L$�@���   �Ѕ��I  �D$�L$���   � UQ�L$�@���   �Ѕ�� U�  �H���   P�D$P�A�С U�L$���@Q�L$�@p�Ѕ���   �D$�L$���   � UQ�L$�@�@|�Ѕ�� U��   �D$�L$���   �@Q�L$�@p�Ѕ���   �D$�L$���   � UQ�L$�@�@p�Ѕ�tl�D$�L$���   � UQ�L$�@�@p�Ѕ�tH�D$�L$���   � UQ�L$�@�@p�Ѕ�t$�D$�L$���   � UQ�L$�@�@p�Ѕ�u� U�@�L$�@��3��@�D$�L$���   � U�@�@�С U�L$Q�@���   �Ѓ��D$    �   � U�L$Q�@�@�Ѓ��3�� U�D$P�I���   �у���_^��]�������̡ UVW���@W�@�С UW�@$�@D�С U�wV�@�@�С UV�@$�@D�Ѓ��G8    �G<   �OH�G@    �GD   �
������S�����������_^��������U���SVW���E�    Q�M��E�    �E�    ������t� �  Q�M��������t� �  Q�M��������t� �  Q�M��������t� �  Q�M�������t� �  Q�M�������t�   Q�M�������t�   Q�M�������t�   Q�M��o�����t� #  Q�M��\�����t� -  Q�M��I�����t� 7  3�9u��~   �]���O��t%� U�U�j R�U��@0�4��@,Q��3ۃ�9]��ËE��W��A��t� Uj SQ�@0R�@�ЋE������W����t� Uj SQ�@0R�@�Ѓ�F;u�|��M���t� UQ�@� �Ѓ�_^[��]���������U��QV��N��t� U�U�j Rh  �@0Q�@,�Ѓ��E����^  �$�`I � Uj j j �@0j j j ���   j h  j<�v�С Uj j j �@0j j j ���   j h  j<�v�С U��P�@0j j j ���   j j j j h"  j<�v�С Uj j j �@0j j j���   j h,  j<�v�Ѓ�Pj j j j j j �  � Uj j j �@0j j j ���   j h  j<�v�С Uj j j �@0j j j ���   j h  j<�v�С U��P�@0j j j ���   j j jj h"  j<�v�С Uj j j �@0j j j���   j h,  j<�v�Ѓ�Pj j j j j j ��  � Uj j j �@0j j j ���   j h  j<�v�С Uj j j �@0j j j���   j h  j<�v�С U��P�@0j j j ���   j j jj h"  j<�v��j j j j j j�  � Uj j j �@0j j j���   j h  j<�v�С Uj j j �@0j j j���   j h  j<�v�С U��P�@0j j j ���   j j jj h"  j<�v��j j j j j j�   � Uj j j �@0j j j���   j h  j<�v�С Uj j j �@0j j j���   j h  j<�v�С U��P�@0j j j ���   j j jj h"  j<�v��j j j j j j � Uj h,  j<�@0�v���   �Ѓ�Pj j j j j j� Uj h6  j<�@0�v���   �Ѓ�(� Uj j j �@0j j j ���   j hy  j�v�С Uj j j �@0j j j ���   j h�  j�v�С U��P�@0j j j ���   j j j j h  j�v�С Uj j j �@0j j j ���   j h  j�v�С U��P�@0j j j ���   j j j j h"  j�v�С Uj j j �@0j j j j ���   h,  j�v�С U��P�@0j j j ���   j j j j h6  j�v�Ѓ�(^��]ÍI �D �E KF �F cG ������������U���  V��W�N��t� U�U�j Rh  �@0Q�@,�Ѓ��N��t� U�U�j Rh  �@0Q�@,�Ѓ��N��t� U�U�j Rh  �@0Q�@,�Ѓ��E�� ��  H��  H�q  �N��t)� Uj j j �@0j j j ���   j h  jQ�Ѓ�(� U������Q�@�@�С U���������@j j�h|7�@Q�ЋN����t.� U������j j j �@0j j j ���   Rh  jQ�Ѓ�(� U������Q�@�@�С U���������@Q�@�С U���������@j j�h�7�@Q�ЋN����t.� U������j j j �@0j j j���   Rh  jQ�Ѓ�(� U������Q�@�@�Ѓ��E�  ���E�    �} �E��jh���h   �tj P�Z�  _^��]� �u�P�I�  _^��]� �N��t)� Uj j j �@0j j j ���   j h  jQ�Ѓ�(� U�M�Q�@�@�С U�M����@j j�h|7�@Q�ЋN����t+� U�U�j j j �@0j j j ���   Rh  jQ�Ѓ�(� U�M�Q�@�@�С U��������@Q�@�С U��������@j j�h�7�@Q�ЋN����t.� U�����j j j �@0j j j���   Rh  jQ�Ѓ�(� U�����Q�@�@�С U�M����@Q�@�С U�M����@j j�h8�@Q�ЋN����t+� U�U�j j j �@0j j j���   Rh  jQ�Ѓ�(� U�M�Q�@�@�Ћ}�E���E�  ���E�    ��jh���h   ���tj ��u�P�j�  �N��t)� Uj j j �@0j j j ���   j h  jQ�Ѓ�(� U������Q�@�@�С U���������@j j�h 8�@Q�ЋN����t.� U������j j j �@0j j j ���   Rh  jQ�Ѓ�(� U������Q�@�@�С U��h������@Q�@�С U��h������@j j�h(8�@Q�ЋN����t.� U��h���j j j �@0j j j���   Rh  jQ�Ѓ�(� U��h���Q�@�@�С U���������@Q�@�С U���������@j j�h08�@Q�ЋN����t.� U������j j j �@0j j jd���   Rh  jQ�Ѓ�(� U������Q�@�@�С U��H������@Q�@�С U��H������@j j�h48�@Q�ЋN����t.� U��H���j j j �@0j j je���   Rh  jQ�Ѓ�(� U��H���Q�@�@�С U�M؃��@Q�@�С U�M؃��@j j�h@8�@Q�ЋN����t+� U�U�j j j �@0j j jf���   Rh  jQ�Ѓ�(� U�M�Q�@�@�С U��(������@Q�@�С U��(������@j j�hD8�@Q�ЋN����t.� U��(���j j j �@0j j jg���   Rh  jQ�Ѓ�(��(���� UQ�@�@�Ѓ��E�  ���E�    �E��jh���h   �����  jP��  _^��]� �N��t)� Uj j j �@0j j j ���   j h  jQ�Ѓ�(� U�M�Q�@�@�С U�Mȃ��@j j�h�7�@Q�ЋN����t+� U�U�j j j �@0j j j���   Rh  jQ�Ѓ�(� U�M�Q�@�@�С U�M����@Q�@�С U�M����@j j�h8�@Q�ЋN����t+� U�U�j j j �@0j j j���   Rh  jQ�Ѓ�(� U�M�Q�@�@�Ћ}�E���E�  ���E�    ��jh���h   ���tj��u�P覱  �N��t)� Uj j j �@0j j j ���   j h  jQ�Ѓ�(� U�M�Q�@�@�С U�M����@j j�h 8�@Q�ЋN����t+� U�U�j j j �@0j j j ���   Rh  jQ�Ѓ�(� U�M�Q�@�@�С U��x������@Q�@�С U��x������@j j�h(8�@Q�ЋN����t.� U��x���j j j �@0j j j���   Rh  jQ�Ѓ�(� U��x���Q�@�@�С U��X������@Q�@�С U��X������@j j�hP8�@Q�ЋN����t1� U��X���j j j �@0j j h�   ���   Rh  jQ�Ѓ�(� U��X���Q�@�@�С U��8������@Q�@�С U��8������@j j�h@8�@Q�ЋN����t1� U��8���j j j �@0j j h�   ���   Rh  jQ�Ѓ�(� U��8���Q�@�@�С U��������@Q�@�С U��������@j j�hT8�@Q�ЋN����t1� U�����j j j �@0j j h�   ���   Rh  jQ�Ѓ�(� U�����Q�@�@�С U���������@Q�@�С U���������@j j�h\8�@Q�ЋN����t1� U������j j j �@0j j h�   ���   Rh  jQ�Ѓ�(� U������Q�@�@�С U���������@Q�@�С U���������@j j�h`8�@Q�ЋN����t1� U������j j j �@0j j h�   ���   Rh  jQ�Ѓ�(� U������Q�@�@�С U���������@Q�@�С U���������@j j�hh8�@Q�ЋN����t1� U������j j j �@0j j h�   ���   Rh  jQ�Ѓ�(� U������Q�@�@�С U���������@Q�@�С U���������@j j�hl8�@Q�ЋN����t1� U������j j j �@0j j h�   ���   Rh  jQ�Ѓ�(� U������Q�@�@�С U��x������@Q�@�С U��x������@j j�ht8�@Q�ЋN����t1� U��x���j j j �@0j j h�   ���   Rh  jQ�Ѓ�(��x��������u�P�O�  _^��]� �������U���<V��N��t*� U�U�j RhM  �@0Q�@,��3���9E������   �N��t*� U�U�j RhN  �@0Q�@,��3���9E������   �N��t*� U�U�j Rh�  �@0Q�@,��3���9E������   �N��t*� U�U�j Rh�  �@0Q�@,��3���9E������   �N��t*� U�U�j Rh  �@0Q�@,��3���9E�����  �N��t*� U�U�j Rh�  �@0Q�@,��3���9E������   �N��t*� U�U�j Rh�  �@0Q�@,��3���9E�����  �N��t*� U�U�j Rh�  �@0Q�@,��3���9E������   �N��t� U�U�j Rh�  �@0Q�@,�Ѓ��N�E���  ��t*� U�U�j Rh�  �@0Q�@,��3���9E������   �N��t*� U�U�j Rh�  �@0Q�@,��3���9E�����  �N��t*� U�U�j Rh�  �@0Q�@,��3���9E������   ��  �E��  P�E��E�    P����  �N��t*� U�U�j Rh�  �@0Q�@,��3���9E������   �N��t� U�U�j Rh�  �@0Q�@,�Ѓ��N�E���,  ��t*� U�U�j Rh  �@0Q�@,��3���9E������   �N��t� U�U�j Rh  �@0Q�@,�Ѓ��N�E���0  ��t*� U�U�j Rh  �@0Q�@,��3���9E������   �N��t� U�U�j Rh  �@0Q�@,�Ѓ��N�E���4  ��t*� U�U�j Rh  �@0Q�@,��3���9E������   �N��t� U�U�j Rh  �@0Q�@,�Ѓ��N�E���8  ��t*� U�U�j Rh#  �@0Q�@,��3���9E������   �N��t� U�U�j Rh%  �@0Q�@0�Ѓ��EȋNfZ���(  ��t*� U�U�j Rh-  �@0Q�@,��3���9E������   �V��t� Uj �H0��$  Ph/  R�A,�Ѓ��N��t*� U�U�j Rh7  �@0Q�@,��3���9E�����   �N��t� U�U�j Rh9  �@0Q�@,�Ѓ��E���<  ^��]���������������U�����E��VW��=�  �A  ��   ����=�   �+  �� ^ �$�^ 3�9�L  ��PQ��D  ��L  ��  ��L  �D$y  �D$�D$    P����  �D$�D$  P���D$    �5�  �   _^��]� 3�9�H  ��PQ��@  ��H  �z�  ��H  �D$�  ��%���j��������   _^��]� ��������   �OX�GH���   �GL���   �GP���   �GT���   P�׹��j �O�-����O��t� UQ�@0�@�Ѓ��� 諰  ������_�   ^��]� �I �\ �] H] v] �]  U������<V���D$DM  ���D$H    �D$Dj jj ���   P軤  ���D$DN  �D$D�D$H    ��j jj ���   P萤  ���D$D�  �D$D�D$H    ��j jj ���   P�e�  ���D$D�  �D$D�D$H    ��j jj ���   P�:�  ���D$D  �D$D�D$H    ��j jj ��  P��  ���D$D�  �D$D�D$H    ��j jj ���   P��  ���D$D�  �D$D�D$H    ��j jj ��  P蹣  �D$8�  ���D$H    j jj ���   �D$T��P莣  ���D$D�  �D$D�D$H    ��jh���h   ���  P�]�  ���D$D�  �D$D�D$H    ��j jj ���   P�2�  ���D$D�  �D$D�D$H    ��j jj ��  P��  ���D$D�  �D$D�D$H    ��j jj ���   P�ܢ  ���D$@�  ��  �D$D    ��P�D$DP�F�  ���D$D�  �D$D�D$H    ��j jj ���   P苢  ���D$D�  �D$D�D$H    jh���h   ���,  P���Z�  ���D$D  �D$D�D$H    ��j jj ���   P�/�  ���D$D  �D$D�D$H    ��jh���h   ���0  P���  ���D$D  �D$D�D$H    ��j jj ���   P�ӡ  ���D$D  �D$D�D$H    ��jh���h   ���4  P袡  ���D$D  �D$D�D$H    ��j jj ���   P�w�  ���D$D  �D$D�D$H    ��jh���h   ���8  P�F�  ���D$D#  �D$D�D$H    ��j jj ���   P��  �D$8%  �D$<    ��<�D$tW���D$,(�:D$��:�D$��(  Z��D$P��  ���D$D-  �D$D�D$H    ��j jj ���   P螠  ���D$D/  �D$D�D$H    ��jh���h   ���$  P�m�  ���D$D7  �D$D�D$H    ��j jj ��   P�B�  ���D$D9  �D$D�D$H    ��jh���h   ���<  P��  ���:����������j �������   ^��]�U����� U��x�@VW���L$�@Q�С U�L$j j�h�6�@Q�@�ЋO����t)� U�T$j j j �@0j j j ���   Rj jQ�Ѓ�(� U�L$Q�@�@�С U�L$Q�@�@�С U�L$ j j�h�6�@Q�@�ЋO����u3��,� U�T$j j j �@0Rj j���   j?h�  Q�Ѓ�$��� U�D$P�I�I�у����?  �O����  � Uj j?h�  �@0Q�@D�Ѓ����w  � U�L$Q�@�@�С U�L$j j�h�6�@Q�@�ЋO����u3��2� U�T$h,  h�  j �@0Rj j���   j?hL  Q�Ѓ�$��� U�D$P�I�I�у�����   � U�L$(Q�@�@�С U�L$,j j�h�6�@Q�@�Ѓ��D$(��P��jhM  辙  � U�L$(Q�@�@�С U�L$,Q�@�@�С U�L$0j j�h�6�@Q�@�Ѓ��D$(��P��jhN  �f�  � U�L$(Q�@�@�ЋO����t� UQ�@0�@X�Ѓ�� U�L$(Q�@�@�С U�L$,j j�h�6�@Q�@�ЋO����u3��2� U�T$(h,  h�  j �@0Rj j���   j?h�  Q�Ѓ�$��� U�D$(P�I�I�у�����   � U�L$Q�@�@�С U�L$j j�h 7�@Q�@�Ѓ��D$��P��jh�  �h�  � U�L$Q�@�@�С U�L$Q�@�@�С U�L$j j�h7�@Q�@�Ѓ��D$��P��jh�  ��  � U�L$Q�@�@�ЋO����t� UQ�@0�@X�Ѓ�� U�L$(Q�@�@�С U�L$,j j�h$7�@Q�@�ЋO����u3��2� U�T$(h,  h�  j �@0Rj j���   j?h  Q�Ѓ�$��� U�D$(P�I�I�у����(  � U�L$Q�@�@�С U�L$j j�h87�@Q�@�Ѓ��D$��P��jh  ��  � U�L$Q�@�@�С U�L$p���@j j��@�С U�L$ljhrab �@�@4�С U�L$Q�@�@�С U�L$j j�hL7�@Q�@�С U�L$���@Qhtitb�L$t�@8�С U�L$Q�@�@�С U�L$p���@jhgbus�@0�С U�L$8Q�@�@�С U�L$<j j�h�6�@Q�@�Ѓ��D$lP���D$HPQhx  ����  ��D  �L$8� UQ�@�@�Ѓ���D   �t  � U�L$HQ�@�@�С U�L$Lj j�hL7�@Q�@�ЋO����u3��,� U�T$Hj j j �@0Rj j���   j9hy  Q�Ѓ�$��� U�D$HP�I�I�у�����  �����g�  Qh�6�L$����j j Q�D$PQjj?h�  ��荒  � U���D$P�I�I�у�����   Qh�6�L$辥���D$��P��jh�  ��  � U�L$Q�@�@��h`7�L$舥��Q�D$��P��h�  ��  � U�L$Q�@�@��h�6�L$�S����D$��P��jh�  �}�  � U�L$Q�@�@�Ѓ���衑  Qh�6�L$����j j Q�D$PQjj?h�  ��藑  � U���D$P�I�I�у����Q  Qh�6�L$�Ȥ���D$��P��jh�  ��  � U�L$Q�@�@��hh7�L$蒤��Q�D$��P��h�  ��  � U�L$Q�@�@�Ѓ���jh�  �
�  Qh|7�L$`�K����D$X�D$�  Pj �D$�D$    P��舑  � U�L$XQ�@�@��h�7�L$`�����D$X�D$�  Pj�D$�D$    P���E�  � U�L$XQ�@�@��h�7�L$`�ţ���D$�  �D$X�D$    Pj�D$��P��  � U�L$XQ�@�@�Ѓ�����  �����  � U�L$Xj j��@�@�С U�L$lj j Q�@�L$d���   �С U�L$X�@�@�С U�L$ljhrab �@�@4�С U�L$HQ�@�@�С U�L$Lj j�h�7�@Q�@�С U�L$\���@Qhtitb�L$t�@8�С U�L$HQ�@�@�С U�L$p���@jhgbus�@0�С U�L$HQ�@�@�С U�L$Lj j�h�6�@Q�@�Ѓ��D$lP���D$XPQh�  ��袍  ��@  �L$H� UQ�@�@�Ѓ���D   �  Qh�7�L$`�+���j j Q�D$dPQjj9h�  ��谎  � U���D$XP�I�I�у�����  �����6�  Qh�6�L$`�ס��j j Q�D$dPQjj?h�  ���\�  � U���D$XP�I�I�у�����   Qh�6�L$`荡���D$X��P��jh�  跐  � U�L$XQ�@�@��h`7�L$`�W���Q�D$\��P��h�  ��  � U�L$XQ�@�@��h�6�L$`�"����D$X��P��j8h�  �L�  � U�L$XQ�@�@�Ѓ����p�  Qh�6�L$`����j j Q�D$dPQjj?h�  ���f�  � U���D$XP�I�I�у���t}Qh�6�L$`蛠���D$X��P��jh�  �ŏ  � U�L$XQ�@�@��h�7�L$`�e���Q�D$\��P��h�  ���  � U�L$XQ�@�@�Ѓ���脎  ��譌  Qh�6�L$`����j j Q�D$dPQjj?h�  ��裌  � U���D$XP�I�I�у����  Qh�6�L$`�ԟ���D$X��P��jh�  ���  � U�L$XQ�@�@��h�7�L$`螟��Q�D$\��P��h�  �)�  � U�L$XQ�@�@�Ѓ���j8h�  ��  Qh�7�L$`�W����D$X�D$�  Pj �D$�D$    P��蔌  � U�L$XQ�@�@��h�7�L$`�����D$X�D$�  Pj�D$�D$    P���Q�  � U�L$XQ�@�@�Ѓ����U�  Qh�6�L$`�ƞ��j j Q�D$dPQjj?h  ���K�  � U���D$XP�I�I�у�����  Qh�6�L$`�|����D$X��P��jh  覍  � U�L$XQ�@�@��h�7�L$`�F���Q�D$\��P��h  �ь  � U�L$XQ�@�@�Ѓ���j8h  辋  Qh�7�L$`������D$X�D$  Pj �D$�D$    P���<�  � U�L$XQ�@�@��h�7�L$`輝���D$X�D$  Pj�D$�D$    P�����  � U�L$XQ�@�@��h�7�L$`�y����D$  �D$X�D$    Pj�D$��P越  � U�L$XQ�@�@��h�7�L$`�6����D$X�D$  Pj�D$�D$    P���s�  � U�L$XQ�@�@��h�7�L$`�����D$X�D$  Pj�D$�D$    P���0�  � U�L$XQ�@�@�Ѓ����4�  Qh�6�L$`襜��j j Q�D$dPQjj?h  ���*�  � U���D$XP�I�I�у�����  Qh�6�L$`�[����D$X��P��jh  腋  � U�L$XQ�@�@��hh7�L$`�%���Q�D$\��P��h  谊  � U�L$XQ�@�@�Ѓ���j8h  蝉  Qh|7�L$`�ޛ���D$X�D$  Pj �D$�D$    P����  � U�L$XQ�@�@��h�7�L$`蛛���D$X�D$  Pj�D$�D$    P���؈  � U�L$XQ�@�@��h�7�L$`�X����D$  �D$X�D$    Pj�D$��P蕈  � U�L$XQ�@�@��h�7�L$`�����D$X�D$  Pj�D$�D$    P���R�  � U�L$XQ�@�@��h8�L$`�Қ���D$X�D$  Pj�D$�D$    P����  � U�L$XQ�@�@�Ѓ�����  Qh�6�L$`脚��j j Q�D$dPQjj?h  ���	�  � U���D$XP�I�I�у����J  Qh�6�L$`�:����D$X��P��jh  �d�  � U�L$XQ�@�@��h8�L$`����Q�D$\��P��h  菈  � U�L$XQ�@�@�Ѓ���j8h  �|�  Qh 8�L$`轙���D$X�D$  Pj �D$�D$    P�����  � U�L$XQ�@�@��h(8�L$`�z����D$X�D$  Pj�D$�D$    P��跆  � U�L$XQ�@�@��h08�L$`�7����D$  �D$X�D$    Pjd�D$��P�t�  � U�L$XQ�@�@��h48�L$`������D$X�D$  Pje�D$�D$    P���1�  � U�L$XQ�@�@��h@8�L$`豘���D$X�D$  Pjf�D$�D$    P����  � U�L$XQ�@�@��hD8�L$`�n����D$X�D$  Pjg�D$�D$    P��諅  � U�L$XQ�@�@��hP8�L$`�+����D$X�D$  Ph�   �D$�D$    P���e�  � U�L$X�@�@Q��h@8�L$`�����D$X�D$  Ph�   �D$�D$    P����  � U�L$XQ�@�@��hT8�L$`蟗���D$X�D$  Ph�   �D$�D$    P���ل  � U�L$XQ�@�@��h\8�L$`�Y����D$X�D$  Ph�   �D$�D$    P��蓄  � U�L$XQ�@�@��h`8�L$`�����D$X�D$  Ph�   �D$�D$    P���M�  � U�L$XQ�@�@��hh8�L$`�͖���D$  �D$X�D$    Ph�   �D$��P��  � U�L$XQ�@�@��hl8�L$`臖���D$X�D$  Ph�   �D$�D$    P�����  � U�L$XQ�@�@��ht8�L$`�A����D$X�D$  Ph�   �D$�D$    P���{�  � U�L$XQ�@�@�Ѓ�����  Qh�6�L$`����j j Q�D$dPQjj?h"  ���u�  � U���D$XP�I�I�у�����   Qh�6�L$`覕���D$X��P��jh#  �Є  � U�L$XQ�@�@��h|8�L$`�p���Q�D$\��P��h$  ���  � U�L$XQ�@�@�Ѓ���h%  �:�  ��賁  Qh�6�L$`�$���j j Q�D$dPQjj?h,  ��詁  � U���D$XP�I�I�у�����   Qh�6�L$`�ڔ���D$X��P��jh-  ��  � U�L$XQ�@�@��h�8�L$`褔��Q�D$\��P��h.  �/�  � U�L$XQ�@�@�Ѓ���h/  �n�  ����  Qh�6�L$`�X���j j Q�D$dPQjj?h6  ���݀  � U���D$XP�I�I�у����  Qh�6�L$`�����D$X��P��jh7  �8�  � U�L$XQ�@�@��h�8�L$`�ؓ��Q�D$\��P��h8  �c�  � U�L$XQ�@�@�Ѓ���j8h9  �P�  Qh�8�L$`葓���D$X�D$9  Pj �D$�D$    P���΀  � U�L$XQ�@�@��h�8�L$`�N����D$X�D$9  Pj�D$�D$    P��苀  � U�L$XQ�@�@�Ѓ����  ���  ���  � U�L$l�@�@�ЋO��t� UQ�@0�@X�Ѓ��O��t� UQ�@0�@X�Ѓ�� U�L$HQ�@�@�С U�L$Lj j�h�8�@Q�@�ЋO����t7� U�T$Rj j �@0�T$Tjj j?Rh�  �D$(    ���   jQ�Ѓ�(� U�L$HQ�@�@�Ѓ��   _^��]á U�L$l�@�@��_3�^��]����������U������4SV���D$     W�L$$�D$Q�u���D$0    �D$4    �  �D$(�\$$���Y  ���؍I � Uh� �@H� �Ћ������  jh�L$ �D$4   �D$<   觍  � Uj ���   �L$4QP�΋B �С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$ QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$Q�Ѓ�� U�L$0Q���   � �С U���΋��   W�@|�С U�L$���   �I�@T�Ћ U��j j �AL�L$�@(�qVR�Ѓ�� Uj �@@�@�Ѓ���K������\$$�D$(��t5�x���x����� UV�@�@�Ѓ���Oy� US�@� �Ѓ�_^[��]� ������������U������$� U�ISV���   �D$    �D$$    W�@4�Ћ����#  ��$    jh�L$���  � Uj ���   �L$$QP�΋B�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$Q�Ѓ�� U�L$ Q���   �@8�Ѓ���uD� U�΋��   �@x��Q�M���w�������t!� UW�I�I�ѡ UWS�@�@�Ѓ�� U�΋��   �@(�Ћ��������� U�L$ Q���   � �Ѓ�_^[��]� ����U������V�uW����   h4  �L$�D$    �D$    茊  � U�L$j QP���   �΋B�ЍL$��  � U�L$Q���   �@H�ЋM��虗������t!� UV�I�I�ѡ UVW�@�@�Ѓ�� U�L$Q���   � �Ѓ�_^��]� �������������������U�� U�� �I���   VW�@T�Ћ U��W�IL�I�ы�����t@�	��$    ��� U�΋��   �@��=�� �  � U�΋��   �@(�Ћ���uˡ Uh�� �@H� �Ћ�������   � U�M�Q�@�@�С U�M�j j�h,9�@Q�@�С U�M������   Q�΋@|�С U�M�Q�@�@�Ѓ��E�   �M��E�@��rje��  � Uj ���   �M�QP�΋B �ЍM��K�  � U�M�Q���   � �С Uj j j �@LVW�@(�Ѓ�� Uj �I@�I�у�_��^��]������U������   SV���D$    W�L$�D$(Q�u���D$     �D$$    �
  �\$3��t$9t$�;  � Uh���@@���   �Ѓ��D$H   �L$<�D$Pn   ��h�  ���  � Uj ���   �L$LQP�ϋB �С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$$Q�L$`Q���   �L$xQR�Ѓ���t(�D$$��t �(U�x`|��t�@`��t
�L$<Q�Ѓ�� U�L$HQ���   � �Ћ���$�   ���D$`   �D$hh�  �-�  � Uj ���   �L$dQP�ϋB �С(U��ub� UjhD �@���   �ЋЃ���tV� U�A�L$ Q�L$HQ���   ��$�   QR�Ѓ���t+�D$ ��t#�(U�x`|��t�@`��t��$�   Q�Ѓ�� U�L$`Q���   � �Ћ U������IRP��$�   P���   �Ћ U������$�   �IP�I�ы U���A��$�   QV�@�С U��$�   Q�@�@�С U��$�   ���@Q�@�С U�L$x���@j j�hD9�@Q�С U�L$<Q�@�@�С U�L$@���@Q�L$xQ�@�С U�L$4���@�@<�Ћ Uj�j��Q��$�   QP�BL�L$<�С U�L$,Q�ϋ��   �@|�С U�L$,Q�@�@�С U�L$x���@Q�@�С U��$�   ���@Q�@�С U���L$(�@Lj W�q��,  �Ћt$��F�t$;t$�������t� US�@� �Ѓ�_^[��]� ��������U������L� USVW�@L�q��(  �Ћ��D$L    ���D$P    �D$8    �D$@    ����  �]�h�  �L$,�r�  � Uj ���   �L$LQP�΋B�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$$QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$(Q�Ѓ�� U�L$HQ���   �@8�Ѓ���n��   h�  �L$4诃  � Uj ���   �L$<QP�΋B�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$$Q���   �L$,QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$0Q�Ѓ�� U�L$8Q���   �@8�Ћˋ�譏����t�8� U�΋��   �@(�Ћ����[���� U�L$8Q���   � �С U�L$LQ���   � �Ѓ�_^[��]� �������U������\S�]VW����  Q�L$4�D$4    �D$8    �D$<    ������t� �  Q�L$4������t� �  Q�L$4������t� �  Q�L$4�ێ����t� �  Q�L$4�ǎ����t� �  Q�L$4賎����t� �  Q�L$4蟎����t� p  Q�L$4苎����t� q  Q�L$4�w�����t� r  Q�L$4�c�����t� s  Q�L$4�O�����t� t  Q�L$4�;�����t� u  Q�L$@�D$@    �D$D    �D$H    ������t� V  Q�L$@�������t� W  Q�L$@������t� X  Q�L$@�Ӎ����t� Y  Q�L$@迍����t� Z  Q�L$@諍����t� [  Q�L$@藍����t� `  Q�L$@胍����t� a  Q�L$@�o�����t� b  Q�L$@�[�����t� c  Q�L$@�G�����t� d  Q�L$@�3�����t� e  �|$4�t$0�L$<�D$X    �D$`    �D$H    �D$P    ���:  �D$0��+��D$���$    �40�L$$�$�  � Uj ���   �L$\QP�ˋB�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$$QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$ Q�Ѓ�� U�L$XQ���   �@8�Ѓ���tW�6�L$,�i  � Uj ���   �L$LQP�ˋB�ЍL$(��~  � U�L$HQ���   �@8�ЋM���֋����t��]�D$��O������t$0� U�L$HQ���   � �С U�L$\Q���   � �ЋL$D����t� UQ�@� �Ѓ���t� UV�@� �Ѓ�_^[��]� �����������U���V���E�   hR  �M��E�   �|~  � U�M�j Q�N���   P�B �ЍM���}  � U�M�Q���   � �Ѓ�^��]���������������U��S�]V3�W9s~$3�� U�U��R�@�@x�Ѕ�t)F��;s|�3�� U�EP�I�I�у���_^[]� �   �������U��M3�V�Q��~�	�u91t@��;�|�3�^]� �   ^]� ��������������U�����U�SWR�E�    �E�    �E�    �P�]3��U�9{~GV�u�3���~���9�t'@;�|���<� ��tQ�M�������t���U�u��EG��;x|�^�E�    _[��t� UR�@� �Ѓ���]� ���U���4��U�SVWR�E�    �E�    �E�    �P�E�E�    �x �3  3ۍI �0�M� U�Q�@�@�С U�M����@QV�@��3���9u�~43����$    �� U�U��M�R�@��@x�Ѕ��!  F��;u�|ء U�M�Q�@�@�С U�MЋ}���@�7Q�@�С U�MЃ��@j j�j �@Q�С U�MЃ��@Q�΋@x�Ћ U����E�P�I�I�у���t7�7Q�M���������t$� UW�I�I�ѡ U���@WV�@�Ѓ��}����EG�}�;x������M���t'�u�Nx!����� U�Q�@�@�ЋM�����Ny��E�    ��t� UQ�@� �Ѓ�_^[��]� � U�M�Q�@�@�Ѓ������������U���VW�}��u����  S�]�d$ � Uj �u�@HW���   �Ѓ�����   ��M�QP���E�    �E�    �E�    �R�}�3�9u�~A�d$ �E3ɋP��~��� 9tA��;�|�EQ���(�����t����}�F;u�|Ƌ]��t� UW�@� �Ѓ��E�    �u��}�E�    �E�    � U�ϋ��   �@4�Ћ��S�uP�R(� U�ϋ��   �@(�Ћ��}������[_^��]� ��������������U���$SV�uW���}�����  �]�d$ � Uj �u�@HV���   �Ѓ����Z  ��M�QP���E�    �E�    �E�    ��u�3��}����   3ɉM�� U�u��M�Q�@�@�С U�M�QV�@�@��3���9s~13���    � U�U܋�R�@�@x�Ѕ��  F��;s|ڋ}� U�M�Q�@�@�ЋE��E��E�6�������t#� UV�I�I�ѡ UV�u�@�@�Ѓ��M�G�u����}�M�;��;����M��tENx'������    � U�Q�@�@�ЋM����Ny��t� UQ�@� �Ѓ��E�    �u�}��E�    �E�    � U�΋��   �@4�Ћ��S�uP�R$� U�΋��   �@(�Ћ��u���H���_^[��]� � U�M�Q�@�@�Ћ}���&������U������(� UVW�q�@L�D$$    �D$,    ��(  �Ћ������
  ��I � U���   �΋R(��h�  �L$���}w  � Uj ���   �L$$QP�΋B�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$Q�Ѓ�� U�L$ Q���   �@8�Ѓ���nu'� U�΋��   �@L�Ѕ�t� UV�@@�@�Ѓ����������� U�L$ Q���   � �Ѓ�_^��]���������������U���   SVW���E�    h�
  �M��E�    �Gv  � U�M���j Q���   �KV�@�ЍM��u  � U�M�Q���   �@8�Ѓ��E�    ���E�    �E�u����E�    P�E�P�  �M���E+��u���@;�L�;�Q�E��P誄���  +����  �	��$    ��� U��l���j hTCAb�@�@�С U��l���h�  hdiem�@�@4�С U��l���jhavem�@�@4�С(U��u[� UjhD �@���   �ЋЃ���tK� U�A�MQ�M�Q���   �M�QR�Ѓ���t&�E��t�(U�x\|��t�@\��t	�M�Q�Ѓ�� U�K�E�    �E�    ���   �@�ЉE��(U�E��
  �E�   ��uW� UjhD �@���   �ЋЃ���tY� U�A�MQ�M�Q���   �M�QR�Ѓ���t4�E��t-�(U�x\|'�ȅ�t!�I\��t�E�P�у��E��M�P�p  �(U��uW� UjhD �@���   �ЋЃ���tQ� U�A�M�Q�M�Q���   �M�QR�Ѓ���t,�E���t%�(U�xx|�ȅ�t�Ix��t�E�P�E�P�у��(U��u[� UjhD �@���   �ЋЃ���tK� U�A�M�Q�M�Q���   �M�QR�Ѓ���t&�EЅ�t�(U�x`|��t�@`��t	�M�Q�Ѓ�� U�K�E�    �E�    �E�    ���   �@T�ЉE܍M��E��E�    �E� UQ�Kj���   �@�С U�M�Q�Kj���   �@�С Uj �@��D  �С(U����u[� UjhD �@���   �ЋЃ���tK� U�A�M�Q�M�Q���   �M�QR�Ѓ���t&�Eԅ�t�(U�x`|��t�@`��t	�M�Q�Ѓ�� U��l����@�@��O�����h�
  �M��r  � Uj ���   �M�Q�KP�B�С(U��u[� UjhD �@���   �ЋЃ���tK� U�A�MQ�MQ���   �M�QR�Ѓ���t&�E��t�(U�x`|��t�@`��t	�M�Q�Ѓ�� U�M�Q���   �@8�Ѓ��E�E��VP�:   �M��t� UQ�@� �Ѓ�� U�M�Q���   � �Ѓ�_^[��]� ����U���,S�]VW3��M��E�    �E�    9;�  ��
  �d$ �F�P�M���p  � Uj ���   �M�QP�E��H�B�С(U��u[� UjhD �@���   �ЋЃ���tK� U�A�MQ�M�Q���   �M�QR�Ѓ���t&�E��t�(U�x`|��t�@`��t	�M�Q�Ѓ�� U�M�Q���   �@�Ѓ���t7� U�M�Q���   �@�Ѓ���u*� U�M�Q���   �@8�Ѓ���uQ�M�|����t�0G��;;������ U�M�Q���   � �Ѓ�_^[��]� ������U��j�h�d�    Pd�%    ��|SVW�e��E�    � U�@�M�Q�@�Ѓ��E�    3��}ܡ U�@�M�@<��;���   � U�@W�MQ�@4������hT9�M��+s���Ћ U�Aj R�@4��f;��á U�@�M�Q�@�Ѓ���tt� U�@W�MQ�@4���� U�@�M�Q�@�Ѓ�� U�@Vj�M�Q�@�Ѓ�� U�@j�j��M�Q�]�S�M̋@L�С U�@�M�Q�@�Ѓ�C�]�G����QhX9�M��rr��Qh\9�M��dr���E�    �E�    � U�@j �M�Q�M�Q�M̋@@�Ѕ���   � U�@j �M�Q�M�Q�M̋@@�Ѕ���   � U�@�M��@<�ЋU�+ЋE�+ЍH� U�@RQ��|���Q�M̋@P�Ћ�� U�I�}W�I�у�� U�AWV�@�С U�@��|���Q�@�Ѓ�� U�@�M�Q�@�Ѓ�� U�@�M�Q�@�Ѓ�� U�H�E�P�I�у�� U�I�EP�I�ы��   �M��y��� U�@�M�Q�@�Ѓ�� U�@�M�Q�@�Ѓ�� U�H�E�P�I�у�� U�I�EP�I���1� U�@�u�@�Ѓ���� ��E������ U�@�MQ�@�ЋE���M�d�    _^[��]� �������U������   SV�u�D$WPV���D$    �D$    �D$    �D$     �D$$    �D$(    �����D$��P�D$P������L$�7x���D$�D$    PV���R����D$��P�D$P������T$��9T$�|$LL$3��L$(���O  �D$�L$h�D$x   Ǆ$�   d   ��HP��k  � Uj ���   �L$|Q�KP�B �С(U��ub� UjhD �@���   �ЋЃ���tS� U�A�L$$Q�L$tQ���   ��$�   QR�Ѓ���t(�D$$��t �(U�x`|��t�@`��t
�L$hQ�Ѓ�� U�L$xQ���   � �С U��$�   ���@Q�@�С U��$�   ���@j j�h\9�@Q�С U��$�   Q�@�@�С U��$�   ���@j j�hX9�@Q�С U�L$@Q�@�@�С U�L$D���@Q��$�   Q�@�С U�L$8���@�@<�Ћ Uj�j�W�Q�L$<P�BL�С U�L$@Q�@�@�С U�L$D���@Q�L$4�@Q�С U�L$H���@�@<�Ћ Uj�j��Q��$�   QP�L$P�BL�С U�L$@�D$P    �D$X    Q���   �L$TQ�@$�С U�L$HQ�@�@�С U�L$<���@Q�@�С U��$�   ���@Q�@�С U��$�   ���@Q�@�ЋD$�L$d���4��i  � Uj ���   �L$TQ�KP�B �С(U��ub� UjhD �@���   �ЋЃ���tS� U�A�L$,Q�L$xQ���   ��$�   QR�Ѓ���t(�D$,��t �(U�x`|��t�@`��t
�L$`Q�Ѓ�� U�L$PQ���   � ��F����;t$(������|$�L$��t� UQ�@� �Ѓ���t<�|$O�\$x!�����I � UV�@�@�Ѓ���Oy� US�@� �Ѓ�_^[��]� U������lSVW���D$H    h�
  �L$$�|$�D$T    �D$\    �D$d    �D$<    �D$D    �h  � U��j ���   �L$LQ�OR�@�ЍL$ �ig  � U�L$H3�Q�t$���   �@8�Ѓ�����  ��
  �C�P�L$,�g  � Uj ���   �L$<Q�OP�B�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$$QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$(Q�Ѓ�� U�L$8Q���   �@�Ѓ����  � U�L$8Q���   �@8�Ѓ���d��   S�L$4��f  � Uj ���   �L$\Q�OP�B�ЍL$0�+f  � U�L$XQ���   �@H�Ћ U������IV�I�ы U���AVW�@�Ѓ��D$xP����� U�L$h�@�@<�Ѕ�t7Q�M�s������t(� UV�I�I�ѡ U�L$l���@VQ�@�Ѓ�� U�L$hQ�@�@�Ћt$���|$� U�L$HF��Q�t$���   �@8�Ѓ�;������ U�L$8Q���   � �С U�L$\�����   Q� �С U�L$L�����   Q� �Ѓ�_^[��]� �U������V�uW����   h�  �L$�D$    �D$    �Le  � U�L$j QP���   �΋B�ЍL$�d  � U�L$Q���   �@H�ЋM���Yr������t!� UV�I�I�ѡ UVW�@�@�Ѓ�� U�L$Q���   � �Ѓ�_^��]� ���U������PVW���D$8   hR  �L$4�D$D   �d  � U�L$8��j Q���   �OV�@ �ЍL$0��c  � U�L$8Q���   � �С U�w�@L��(  �Ѓ��D$H    �D$P    ������  �(U��ut� UjhD �@���   �ЋЃ�����   � U�A�L$Q�L$Q���   �L$$QR�Ѓ�����   �L$����   �(U�y\��   ����   �A\����   �L$0Q�С(U���D$8�  �D$<    �D$@    ��u_� UjhD �@���   �ЋЃ���tU� U�A�L$Q�L$$Q���   �L$,QR�Ѓ���t-�D$��t%�(U�xd|��t�@d��t�L$8Q�L$4Q�Ѓ�� U�L$Hj Q�L$8���   Q�΋@�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$,Q���   �L$4QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$0Q�Ѓ�� U�L$HQ���   �@8�Ѓ�����   � U�΋��   �@(�������� Uh���@@���   �Ѓ��D$8   �L$0�D$@   ��h�  ��a  � Uj ���   �L$<QP�΋B �ЍL$0�Va  � U�L$8Q���   � �С Uj V�w�@L��,  �Ѓ�� U�L$HQ���   � �Ѓ�_^��]������������̡ UV�q�@L���   �Ћ U�������   �΋R��=�� t+� U�΋��   �@(�С U�΋��   �@��=�� uՋ�^�������������������������������U������4S��VW�{ �.  �D$$�D$$    P�u�D$0    �D$4    �3����|$(3�����   ��I �D$$�L$��R  P�`  � U�L$0�D$0   �D$8   j ���   Q�L$$Q�K�@ �С U�L$0Q���   � �С(U����u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$ QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$Q�Ѓ�F;��"����L$$��t� UQ�@� �Ѓ�_^[��]� �U������,S�]V�   �L$W�D$(    �D$0    �~��I ��R  P�L$$�p_  � U�L$(j Q�L$(���   Q�L$�@�I�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$$QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$ Q�Ѓ�� U�L$(Q���   �@�Ѓ���u*� U�L$(Q���   �@8�Ѓ���tQ���Ck����t�0FO����� U�L$(Q���   � �Ѓ�_^[��]� �����U������V�u����   h  �L$�D$    �D$    �-^  � U�L$j QP���   �΋B�ЍL$�]  � U�L$Q���   �@8��H����w%� U�L$Q���   �@8�ЋM���|j����t�0� U�L$Q���   � �Ѓ�^��]� ��������U������PVW��� t]h�  �L$4�]  � U�L$8�D$8   �D$@   j ���   Q�L$8Q�O�@ �С U�L$8Q���   � �Ѓ��L$0�\  � t]h  �L$4�]  � U�L$8�D$8   �D$@   j ���   Q�L$8Q�O�@ �С U�L$8Q���   � �Ѓ��L$0�M\  hR  �L$4�D$<   �D$D   �\  � U��j ���   �L$<Q�OR�@ �ЍL$0�\  � U�L$8Q���   � �С U�w�@L��(  �Ѓ��D$H    �D$P    ������  �(U��ut� UjhD �@���   �ЋЃ�����   � U�A�L$Q�L$Q���   �L$$QR�Ѓ�����   �L$����   �(U�y\��   ����   �A\����   �L$0Q�С(U���D$8�  �D$<    �D$@    ��u_� UjhD �@���   �ЋЃ���tU� U�A�L$Q�L$$Q���   �L$,QR�Ѓ���t-�D$��t%�(U�xd|��t�@d��t�L$8Q�L$4Q�Ѓ�� U�L$Hj Q�L$8���   Q�΋@�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$,Q���   �L$4QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$0Q�Ѓ�� U�L$HQ���   �@8�Ѓ�����   � U�΋��   �@(�������� Uh���@@���   �Ѓ��D$8   �L$0�D$@   ��h�  �Z  � Uj ���   �L$<QP�΋B �ЍL$0�pY  � U�L$8Q���   � �С Uj V�w�@L��,  �Ѓ�� U�L$HQ���   � �Ѓ�_^��]�������U���(VW��3��d$ ��S  P�M��Y  � U�M��E�   �E�    j ���   Q�M�Q�O�@ �С U�M�Q���   � �С(U����u[� UjhD �@���   �ЋЃ���tK� U�A�M�Q�M�Q���   �M�QR�Ѓ���t&�E���t�(U�x`|��t�@`��t	�M�Q�Ѓ�F���2���_^��]������������̡ UV�q�@L���   �Ћ U�������   �΋R��=�� t+� U�΋��   �@(�С U�΋��   �@��=�� uՋ�^���������������U������D  SVW�D$�D$    P�u���D$$    �D$(    �z����L$�VUUU������t$0�v+�tF�t$0h  �L$(Ǆ$�       Ǆ$�       ��W  � U��j ���   ��$�   Q�OR�@�ЍL$$�W  � U��$�   Q���   �@8�й@   Ǆ$4      +�Ǆ$<      ���L$t3�;Ή\$,��L�;ء U���   �^  �@8��$�   Q�Ѓ�Ǆ$h     ��$�  �p�h  ��$t  �W  � Uj ���   ��$l  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$HQ��$�  Q���   ��$�  QR�Ѓ���t+�D$H��t#�(U�x`|��t�@`��t��$�  Q�Ѓ�� U��$h  Q���   � �С U���@j ��D  �Ѝ�  �D$�� �D$���(U�D$    Ǆ$�     Ǆ$�     Ǆ$�   �  Ǆ$�       Ǆ$�       ��ue� UjhD �@���   �ЋЃ���tu� U�A�L$PQ��$�  Q���   ��$  QR�Ѓ���tG�D$P��t?�(U�x\|4��t0�@\��t)�L$<Q�Ѓ��D$�L$<P��Q  ��$�   P�L$@�7Q  � U��$�  j Q�L$D���   Q�O�@ �С(U��uk� UjhD �@���   �ЋЃ���t\� U�A��$�   Q��$X  Q���   ��$l  QR�Ѓ���t+��$�   ��t �(U�x`|��t�@`��t
�L$<Q�Ѓ�� U��$�  Q���   � �С(U��Ǆ$�     Ǆ$�     Ǆ$�   �  Ǆ$�       Ǆ$�       ��ue� UjhD �@���   �ЋЃ���tu� U�A�L$DQ��$  Q���   ��$�  QR�Ѓ���tG�D$D��t?�(U�x\|4��t0�@\��t)�L$4Q�Ѓ��D$�L$4P�BP  ��$�   P�L$8�O  � U��$�  j Q�L$<���   Q�O�@ �С(U��uk� UjhD �@���   �ЋЃ���t\� U�A��$�   Q��$�  Q���   ��$�  QR�Ѓ���t+��$�   ��t �(U�x`|��t�@`��t
�L$4Q�Ѓ�� U��$�  Q���   � �Ѝ[���p�X;D$�  �L$����$  ��$�  ��$|  P�D$Ǆ$�     PǄ$�  �  Ǆ$�      Ǆ$�      �O  � Uj ���   ��$�  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$|Q��$�  Q���   ��$�  QR�Ѓ���t+�D$|��t#�(U�x`|��t�@`��t��$  Q�Ѓ�� U��$�  Q���   � �Ѓ��D$;��  �D$��$�  ����$�  ��$�   P�D$Ǆ$�     PǄ$�   �  Ǆ$�       Ǆ$�       �N  � Uj ���   ��$�  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$LQ��$�  Q���   ��$�  QR�Ѓ���t+�D$L��t#�(U�x`|��t�@`��t��$�  Q�Ѓ�� U��$�  Q���   � �ЋD$ ��;��  �D$��$  ����$�  ��$@  P�D$Ǆ$�     PǄ$H  �  Ǆ$L      Ǆ$P      �M  � Uj ���   ��$�  Q�OP�B �С(U��uk� UjhD �@���   �ЋЃ���t_� U�A��$�   Q��$�  Q���   ��$�  QR�Ѓ���t.��$�   ��t#�(U�x`|��t�@`��t��$  Q�Ѓ�� U��$�  Q���   � �Ѓ�� U�\$,�H�ÙRP��$H  P���   �Ћ U������$�  �IP�I�ы U���A��$�  QV�@�С U��$H  Q�@�@�С U��$  ��Ǆ$�      Ǆ$�      ���   Q��$�  Q�@$�С(U��Ǆ$�   �  Ǆ$�       Ǆ$       ��ue� UjhD �@���   �ЋЃ���tu� U�A�L$TQ��$�  Q���   ��$   QR�Ѓ���tG�D$T��t?�(U�x\|4��t0�@\��t)�L$$Q�Ѓ��D$�L$$P��J  ��$�   P�L$(�J  � U��$�  j Q�L$,���   Q�O�@ �С(U��uk� UjhD �@���   �ЋЃ���t\� U�A��$�   Q��$  Q���   ��$  QR�Ѓ���t+��$�   ��t �(U�x`|��t�@`��t
�L$$Q�Ѓ�� U��$�  Q���   � �С U��$�  ���@Q�@�Ѓ�� ��   ��$p  Ǆ$     P�D$Ǆ$     P��$  Ǆ$x  �  Ǆ$|      Ǆ$�      �,J  � Uj ���   ��$  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$`Q��$  Q���   ��$,  QR�Ѓ���t+�D$`��t#�(U�x`|��t�@`��t��$  Q�Ѓ���$  ��   �GL��$  ��$0  ��$  P�D$Ǆ$,     PǄ$  �  Ǆ$      Ǆ$       �0I  � Uj ���   ��$,  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$\Q��$4  Q���   ��$D  QR�Ѓ���t+�D$\��t#�(U�x`|��t�@`��t��$  Q�Ѓ���$(  � UQ���   � �Ѓ��  �  �GP��$�  ��$H  ��$X  P�D$Ǆ$D     PǄ$`  �  Ǆ$d      Ǆ$h      �H  � Uj ���   ��$D  Q�OP�B �С(U��uk� UjhD �@���   �ЋЃ���t_� U�A��$�   Q��$L  Q���   ��$\  QR�Ѓ���t.��$�   ��t#�(U�x`|��t�@`��t��$�  Q�Ѓ�� U��$@  Q���   � �Ѓ��$ �
  �GT��$(  ��$`  ��$(  P�D$Ǆ$\     PǄ$0  �  Ǆ$4      Ǆ$8      �G  � Uj ���   ��$\  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$hQ��$d  Q���   ��$�  QR�Ѓ���t+�D$h��t#�(U�x`|��t�@`��t��$(  Q�Ѓ�� U��$X  Q���   � �Ѓ��( �}  � U��$l  Q�@�@�С U���H��$l  P�GXP�A�С U��$t  Ǆ$�      Ǆ$�      Q���   ��$�  Q�@$�Ѓ�Ǆ$�   p  ��$�   Ǆ$�       ��$   Ǆ$�       P�D$P�E  � Uj ���   ��$�  Q�OP�B �С(U��uk� UjhD �@���   �ЋЃ���t_� U�A��$�   Q��$�  Q���   ��$p  QR�Ѓ���t.��$�   ��t#�(U�x`|��t�@`��t��$   Q�Ѓ�� U��$�  Q���   � �С U��$p  ���@Q�@�Ѓ��4 �
  �Gp��$4  ��$�  ��$�   P�D$Ǆ$�     PǄ$�   q  Ǆ$�       Ǆ$�       �gD  � Uj ���   ��$�  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$pQ��$�  Q���   ��$�  QR�Ѓ���t+�D$p��t#�(U�x`|��t�@`��t��$4  Q�Ѓ�� U��$�  Q���   � �Ѓ��8 �  �Gt��$$  ��$�  ��$�   P�D$Ǆ$�     PǄ$�   r  Ǆ$�       Ǆ$�       �SC  � Uj ���   ��$�  Q�OP�B �С(U��uk� UjhD �@���   �ЋЃ���t_� U�A��$�   Q��$�  Q���   ��$�  QR�Ѓ���t.��$�   ��t#�(U�x`|��t�@`��t��$$  Q�Ѓ�� U��$�  Q���   � �Ѓ��< �
  �Gx��$@  ��$�  ��$  P�D$Ǆ$�     PǄ$  s  Ǆ$      Ǆ$      �9B  � Uj ���   ��$�  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$xQ��$�  Q���   ��$�  QR�Ѓ���t+�D$x��t#�(U�x`|��t�@`��t��$@  Q�Ѓ�� U��$�  Q���   � �Ѓ��@ �  �G|��$8  ��$�  ��$  P�D$Ǆ$�     PǄ$$  t  Ǆ$(      Ǆ$,      �%A  � Uj ���   ��$�  Q�OP�B �С(U��uk� UjhD �@���   �ЋЃ���t_� U�A��$�   Q��$�  Q���   ��$�  QR�Ѓ���t.��$�   ��t#�(U�x`|��t�@`��t��$8  Q�Ѓ�� U��$�  Q���   � �Ѓ��0 �  �Gl��$4  Z�P�D$Ǆ$�     P��$T  Ǆ$<  w  Ǆ$@      Ǆ$D      ��$�  �@  � Uj ���   ��$�  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$XQ��$�  Q���   ��$�  QR�Ѓ���t+�D$X��t#�(U�x`|��t�@`��t��$L  Q�Ѓ�� U��$�  Q���   � �Ѓ��, �
  �Gh��$�  ��$   ��$L  P�D$Ǆ$�     PǄ$T  v  Ǆ$X      Ǆ$\      ��>  � Uj ���   ��$�  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$dQ��$�  Q���   ��$4  QR�Ѓ���t+�D$d��t#�(U�x`|��t�@`��t��$�  Q�Ѓ�� U��$�  Q���   � �Ѓ��D �  ���   ��$X  ��$  ��$d  P�D$Ǆ$     PǄ$l  u  Ǆ$p      Ǆ$t      ��=  � Uj ���   ��$  Q�OP�B �С(U��ue� UjhD �@���   �ЋЃ���tY� U�A�L$lQ��$�  Q���   ��$�  QR�Ѓ���t+�D$l��t#�(U�x`|��t�@`��t��$X  Q�Ѓ�� U��$  Q���   � �Ѓ��t$0C�L$t����� ��$0  Q�С U��$�   �����   Q� �ЋL$����t� UQ�@� �Ѓ�_^[��]� ������U������  SVW��Ǆ$�       h�  �L$T�\$Ǆ$�       �W?  � U��$�   ��j Q���   �KV�@�ЍL$P�>  � U��$�   Q���   �@8�Ѓ����  h  ��$�   �D$4    �D$<    ��>  � Uj ���   �L$4Q�KP�B�Ѝ�$�   �@>  � U�L$0Ǆ$      3�Ǆ$      Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       �D$X    �D$`    �D$@    �D$H    �D$     �D$(    ���   Q�@8�Ѓ�����  �}���$    ��  �D$�� �D$��$�   �D$l�D$    P�D$�D$p�  P�D$x    �D$|    �;  � Uj ���   ��$�   Q�KP�B�С(U��ub� UjhD �@���   �ЋЃ���tV� U�A�L$Q��$�   Q���   �L$XQR�Ѓ���t+�D$��t#�(U�x`|��t�@`��t��$�   Q�Ѓ�� U��$�   Q���   �@8�Ѓ����m  ��$�   Ǆ$�   �  P�D$Ǆ$�       P��$�   Ǆ$�       �:  � Uj ���   ��$�   Q�KP�B�Ѝ�$�   �1<  � U��$�   Q���   �@8�Ѓ�����  ��$�   Ǆ$�   �  P�D$Ǆ$�       P��$  Ǆ$�       �9  � Uj ���   �L$\Q�KP�B�Ѝ�$  �;  �D$x�D$x�  P�D$Ǆ$�       P��$   Ǆ$�       �'9  � Uj ���   �L$DQ�KP�B�Ѝ�$�   �O;  ��$�   Ǆ$�   �  P�D$Ǆ$�       P��$  Ǆ$�       ��8  � Uj ���   �L$$Q�KP�B�Ѝ�$   ��:  � U�L$XQ���   �@8�Ѓ���t$� U�L$XQ���   �@8�Ћϋ���G����t�� U�L$@Q���   �@8�Ѓ���t$� U�L$@Q���   �@8�Ћϋ��G����t�� U�L$ Q���   �@8�Ѓ���t$� U�L$ Q���   �@8�Ћϋ��cG����t��\$� U�L$0QF���   �@8�Ѓ�;��h���� U�L$ Q���   � �С U�L$DQ���   � �С U�L$`Q���   � �С U��$�   Q���   � �С U��$�   Q���   � �С U��$$  Q���   � �С U�L$HQ���   � �Ѓ�� U��$�   Q���   � �Ѓ�_^[��]� �������������U������V�u����   h�  �L$�D$    �D$    �9  � Uj ���   �L$QP�΋B�ЍL$��8  � U�L$Q���   �@8�Ѓ���tsh�  �L$�?9  � U�L$j QP���   �΋B�ЍL$�8  � U�L$Q���   �@8�Ѓ���t%� U�L$Q���   �@8�ЋM���E����t�0� U�L$Q���   � �Ѓ�^��]� ������������U������PVW���D$8   hR  �L$4�D$D   �8  � U�L$8��j Q���   �OV�@ �ЍL$0��7  � U�L$8Q���   � �С U�w�@L��(  �Ѓ��D$H    �D$P    ������  �(U��ut� UjhD �@���   �ЋЃ�����   � U�A�L$Q�L$Q���   �L$$QR�Ѓ�����   �L$����   �(U�y\��   ����   �A\����   �L$0Q�С(U���D$8�  �D$<    �D$@    ��u_� UjhD �@���   �ЋЃ���tU� U�A�L$Q�L$$Q���   �L$,QR�Ѓ���t-�D$��t%�(U�xd|��t�@d��t�L$8Q�L$4Q�Ѓ�� U�L$Hj Q�L$8���   Q�΋@�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$,Q���   �L$4QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$0Q�Ѓ�� U�L$HQ���   �@8�Ѓ�����   � U�΋��   �@(�������� Uh���@@���   �Ѓ��D$8   �L$0�D$@   ��h�  ��5  � Uj ���   �L$<QP�΋B �ЍL$0�F5  � U�L$8Q���   � �С Uj V�w�@L��,  �Ѓ��D$8   �L$0�D$@   h�  �{5  � Uj ���   �L$<Q�OP�B �ЍL$0��4  � U�L$8Q���   � �Ѓ�� U�L$HQ���   � �Ѓ�_^��]��̡ UV�q�@L���   �Ћ U�������   �΋R��=�� t+� U�΋��   �@(�С U�΋��   �@��=�� uՋ�^���������������U������  SVW�D$�D$    P�u���D$    �D$     ����3��|$9|$�^  ���$    �� Uh�� �@H� �Ћ�����u� UV�@@�@���  �D$� U���I�D$$� �RP��$   P���   �Ћ U������$�   �IP�I�ы U���A��$�   QW�@�С U��$   Q�@�@�С U��$�   ���@Q�@�С U�L$|���@j j�hd9�@Q�С U�L$lQ�@�@�С U�L$p���@Q�L$|Q�@�С U�L$d���@�@<�Ћ Uj�j��Q��$�   QP�L$l�BL�С U�L$\Q�΋��   �@|�С U�L$\Q�@�@�С U�L$|���@Q�@�С U��$�   ���@Q�@�Ѓ��L$4h�  ��2  � U��$�   Ǆ$�      Ǆ$�   |  j ���   Q�L$<Q�@ ���С U��$�   Q���   � �С(U����ub� UjhD �@���   �ЋЃ���tS� U�A�L$(Q�L$xQ���   ��$�   QR�Ѓ���t(�D$(��t �(U�x`|��t�@`��t
�L$4Q�Ѓ�h  �L$H��1  �L$$j ���$�   ��$�   � UǄ$�      Q�L$L���   Q�΋@ �С U��$�   Q���   � �С(U����ue� UjhD �@���   �ЋЃ���tV� U�A�L$0Q��$   Q���   ��$�   QR�Ѓ���t(�D$0��t �(U�x`|��t�@`��t
�L$DQ�Ѓ�hx  �L$X�	1  �C��$�   ��$�   � UǄ$�      j Q���   �L$\Q�΋@ �С U��$�   Q���   � �С(U����ue� UjhD �@���   �ЋЃ���tV� U�A�L$,Q��$�   Q���   ��$�   QR�Ѓ���t(�D$,��t �(U�x`|��t�@`��t
�L$TQ�Ѓ�h�  �L$@�,0  �C��$�   ��$�   � UǄ$�      j Q���   �L$DQ�΋@ �С U��$�   Q���   � �С(U����ub� UjhD �@���   �ЋЃ���tS� U�A�L$ Q��$  Q���   �L$xQR�Ѓ���t(�D$ ��t �(U�x`|��t�@`��t
�L$<Q�Ѓ�h  �L$P�R/  � U��$   Ǆ$      Ǆ$     j ���   Q�L$TQ�@ ���С U��$   Q���   � �С(U����ub� UjhD �@���   �ЋЃ���tS� U�A�L$Q�L$pQ���   ��$�   QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$LQ�Ѓ�� U�K ���   �@x�Ћ UP�A�@�С U���K���   �@T�Ћ U��j j �s �ALVR�@(�С U���@@j �@�Ћ|$G���|$;|$������L$��t� UQ�@� �Ѓ�_^[��]� �����������U������L� U�I SV���   W�@4�Ћ��D$H    �D$P    �D$8    �D$@    ����  �]�d$ h�  �L$,�-  � U�L$Hj Q�L$0���   Q�΋@�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$Q���   �L$$QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$(Q�Ѓ�� U�L$HQ���   �@8�Ѓ�=|  ��   h  �L$4�,  � U�L$8j Q�L$8���   Q�΋@�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$$Q���   �L$,QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$0Q�Ѓ�� U�L$8Q���   �@8�Ѓ���t$� U�L$8Q���   �@8�Ћˋ��8����t�8� U�΋��   �@(�Ћ����7���� U�L$8Q���   � �С U�L$LQ���   � �Ѓ�_^[��]� ���U������V�u��t~hw  �L$�D$    �D$    �a+  � U�L$j QP���   �΋B�ЍL$�*  � U�L$Q���   �@8�ЋM����7����t�0� U�L$Q���   � �Ѓ�^��]� ����������U������PVW���D$8   hR  �L$4�D$D   ��*  � U�L$8��j Q���   �OV�@ �ЍL$0�*  � U�L$8Q���   � �С U�w�@L��(  �Ѓ��D$H    �D$P    ������  �(U��ut� UjhD �@���   �ЋЃ�����   � U�A�L$Q�L$Q���   �L$$QR�Ѓ�����   �L$����   �(U�y\��   ����   �A\����   �L$0Q�С(U���D$8�  �D$<    �D$@    ��u_� UjhD �@���   �ЋЃ���tU� U�A�L$Q�L$$Q���   �L$,QR�Ѓ���t-�D$��t%�(U�xd|��t�@d��t�L$8Q�L$4Q�Ѓ�� U�L$Hj Q�L$8���   Q�΋@�С(U��u_� UjhD �@���   �ЋЃ���tP� U�A�L$Q�L$,Q���   �L$4QR�Ѓ���t(�D$��t �(U�x`|��t�@`��t
�L$0Q�Ѓ�� U�L$HQ���   �@8�Ѓ�����   � U�΋��   �@(�������� Uh���@@���   �Ѓ��D$8   �L$0�D$@   ��h�  �*(  � Uj ���   �L$<QP�΋B �ЍL$0�'  � U�L$8Q���   � �С Uj V�w�@L��,  �Ѓ�� U�L$HQ���   � �Ѓ�_^��]�������������U���(� U�I VW���   �@8�Ћ��E�    �E�    ���  ���$    �d$ � U�����   �ϋ@,��h�  �M���L'  � U�M�j Q�M싀�   Q�΋@�С(U��u[� UjhD �@���   �ЋЃ���tK� U�A�M�Q�M�Q���   �M�QR�Ѓ���t&�E���t�(U�x`|��t�@`��t	�M�Q�Ѓ�� U�M�Q���   �@8�Ѓ�=|  u'� U�΋��   �@L�Ѕ�t� UV�@@�@�Ѓ��������� U�M�Q���   � �Ѓ�_^��]����U��q �s8  � U�IV���   �@T�Ћ U��h�� R�AL���   �Ћȃ���u3�^��]á U�� ���j h'  R���   ���   ������������������ U���   �@X�Ћȅ�u"��� ��'  � U����   �@X�Ћȅ�t�� U���   �@(�Ћ U�Ћ��   �ʋ@(�Ћ U�Ћ��   �ʋ@(��^��]��������������̡ UV�q�@L���   �Ћ U�������   �΋R��=�� t+� U�΋��   �@(�С U�΋��   �@��=�� uՋ�^����������������k  �����������U��=dU �hU   ui� UVh�9jU�@j���   �Ћ�����t3� UV�I�I�ѡ UV�@$�@D�С UV�u�@$�@L�Ѓ��3��5dU��^u3�]� �=\U t3�9XU��]� � U�u�@<� �Ћ��\U   3��XU������]� ����������U�������   S3�VW����$�   98UtC�L$,�   � +  ���L$H�D$P� *  ���Y)  � U��VR�A$�@<�Ѓ��D$��u�D$ ��t-� U�L$Q����@$�@H�С U�L$���@Q�@�Ѓ���t-� U�L$HQ����@$�@H�С U�L$L���@Q�@�Ѓ���t*� U�L$,Q�@$�@H�С U�L$0���@Q�@�Ѓ��|$ � U�@�@��  �58U��$�   Q�С U��$�   ���@$Q�@D�С U��$�   ���@$QV�@L�С U��$�   Q�@$�@h�Ѓ���$�   ��$�   P�'  � U���D$P�I�I�ы U���A$�L$Q�@D�С U�L$���@$VQ�@�С U�L$PQ�@�@�С U�L$T���@$Q�@D�С U�L$L���@$hp9Q�@d�С U�L$4Q�@�@�С U���@$�L$,Q�@D�С U�L$0���@$hx9Q�@d�Ѝ�$�   �)  � U���D$lP�I�I�ы U���A$�L$dQ�@D�С U�L$h���@$QV�@L�С U�L$4Q�L$pQ�@$�@@�С U��$�   Q�@�@�С U��$�   ���@$Q�@D�С U��$�   ���@$Q�L$hQ�@L�С U�L$PQ��$�   Q�@$�@@�С UW�@�@�Ѓ�� UW�@$�@D�С U��$�   ���@$WQ�@L�С U�L$QW�@$�@@�С U��$�   Q�@$�@H�С U��$�   ���@Q�@�С U�L$h���@$Q�@H�С U�L$h���@Q�@�С U��$�   ���@$Q�@H�С U��$�   ���@Q�@�С U�L$0���@$Q�@H�С U�L$0���@Q�@�С U�L$L���@$Q�@H�С U�L$L���@Q�@�С U�L$���@$Q�@H�С U�L$���@Q�@�С U��$�   ���@Q�@�С U��$�   ���@$Q�@H�Ѝ�$�   ��   �L$Q�С U�L$���@$Q�@D�С U�L$���@$h�9Q�@d�Ѝ�$�   �%  � U��W�I�I�ы U���A$W�@D�С U���@$WV�@L�С U�L$QW�@$�@@�С U��$�   Q�@$�@H�С U��$�   ���@Q�@�С U�L$���@$Q�@H�ЍL$� U���@Q�@�Ѓ���_^[��]������������̃=`U uz�XU��t!� U�5hUQ�@<�@�Ѓ��XU    V�5dU��tC� UV�@$�@H�С UV�@�@�ЋdU����t� UQ�@� �Ѓ��dU    ^��������������k���������������XU    �XU�\U    �dU    �`U    ���U���VQ�M�����P����� U���E�P�I$�IH�ы U�A�M�Q�@�Ѓ���^��]����������̋� U��������V���t�j �� UV�@� �Ѓ�^����9������������9����������U���u�M�u�u��u�P]��������U��M�u�u��P]��������������U��M�u��P]�U��M�]� ����̡ UQ�@L���   �Ѓ�������������U�� Uj �u�@LQ��,  �Ѓ�]� � UQ�@L��(  �Ѓ�������������U�� Uj j �u�@L�uQ�@(�Ѓ�]� �������������̡ UQ�@L�@,�Ѓ���������������̡ UQ�@L�@�Ѓ���������������̸   � ��������U�� U�u�H�I�ыE��]� ��̸   � ��������3�� ����������̸   @� ��������3�� �����������3�� ����������̸   � ��������U����   V�uW����u3�_^��]�h�   ��@���j P�s-  �E��@����E�� Uh�   QW�@h� ��`����E�    ǅ@���   ǅD���@� �E�] �E�S �E�l �E�X �E�v �E�b �E�g �E�q ���   jh�>  �Ѓ�$_^��]ËI �$U    ��t� UjQ�@P�@�Ѓ�� Uj�@�@,�Ѓ�3������������������������̋A��uË ����̋A�������������U��V���PD��t�E9Ft
�F�΋�PH^]� ����������U���� UV�u�V�E�    �    �B    ��������   �E�j P�E�    �IR�ы U�E�P���   �	�у���^��]� �����������3�� �����������3���������������3���������������3�������������������������������3���������������3���������������U�� UV��M�@�@ ��=ytsdt�u���u�6   ^]� � U�v�@0���   �Ћ�����P�   ^]� ����������U�� UV��M�@�@ ��=cksat]=ckhct�u���u�?  ^]� � Uj j j j j j j �F   �@0j j �v���   �Ѓ�(��t#�F    �   ^]� �~ t����P^]� 3�^]� �������������V��N��9��t� UQ�@0�@�Ѓ��F    ^�������U��Q� USVW�@�ً}3��ω]��@ ��=INIb�  ��   =SACbmt)=$'  t
=MicM�}  ���W�P$�   _��^[��]� ��MQ�M��u�Q�ˉu�P��t� U�u�u��@4�s�@�Ѓ��   _��^[��]� =ARDb�  � U��j j�@���   �Ћ؋ϡ Uj j�@���   �ЋM��� Uj j�@���   �ЋM�� Uj j�@���   ���u�M�PVW�S�R�   _��^[��]� ����P�   _��^[��]� =NIVbvt]=NPIbtE=ISIbum� U�s�@4�@���s�� U�@4�@�Ћ����VP�R�   _��^[��]� ���W�P_^[��]� ����P�   _��^[��]� =cnyst_��^[��]� � U��j hIicM�@���   �Ћ��WP�R _^[��]� � �������������3�� ������������ �������������3�� ����������̸   � ��������U���u��u�u�u�P]� ��������U�� UV��h�  �@4�v�@$���u� U�u�u�@4�u�v�@�Ѓ�2�^]� ��������������̸   ����������̸   ����������̡ Uh�  �q�@4�@$�Ѓ�� �����U���u� U�u�u�@4�u�q�@�Ѓ�]� ���������̡ U�q�@4�@�Ѓ�������������̡ U�q�@4�@�Ѓ��������������V��~ �:u� U�v�@4� �Ѓ��F    �F    ^����������������U�� US�]V�@��ˋ@ ��=ckhc��   t|=cksatb=TCAb��   � U��Wj hdiem�@���   �Ћ��SW���F   �R�~ ��t��t��u3��΃���P�   _^��[]� �~ ti����P^[]� �~ tV� Uj j j �@0j j j ���   j j j �v�Ѓ�(��t*�F    �   ^[]� =atnit�u��S��  ^[]� ^3�[]� ����������U��E�A�I��u3�]� � UQ�@0�@�Ѓ�]� �����V��N��9��t� UQ�@0�@�Ѓ��F    ^�������3�� ����������̸   ����������̡ Uj j j �@0j j j ���   j j j �q�Ѓ�(��������U���V�q��u�E�    �p^��]� �E�H�� UQ�u�M�@0RVQ���   �Ћu� Uj P�    �F    ���   V�I�ы U�E�P���   �	�у�$��^��]� �������̡ U�q�@0���   �Ѓ�����������U�� U�M���@Vj j��@�ЋM� U��t �@4Q�@�Ѓ���t$��M�Q�u���R(�$�@0�u�@�Ћȃ���u3��:��U�R�u�P ���M� U�@�@ �Ѓ��t� U�M�Q�u�@0�@x�Ѓ�� U�Q�M�R�ҋ�^��]�����������������$U    ������U���� UV�u ��M�@j��@�С U�M�h/D h8kds�@�@4�С U�M Q�M��E     Q�@0j jj ���   j9�u�uj2�v�Ћ U��(�u �Q�M�R�ҋ�^��]� ������U��EV�P�0� URj j �@0j j �u���   j Vj<�q�Ѓ�(^]� ��������U��Ej j j �� Uj j j �@0j Rj�q���   �Ѓ�(]� ������������̋I��u3�� � Uj j
j �@0j
Q�@T�Ѓ�� �������̋I��u3�á UQ�@0�@X�Ѓ������U��I��u3�]�  �u$� U�u j �u�@0j �u�u���   �uQ�Ѓ�$]�  �̋I��u3�� � Uj j?h�  �@0Q�@D�Ѓ�� �������U��V�q��u3�^]� �E�H�� UQj j �@0j j j ���   j RjV�Ѓ�(^]� �������������U��V�q��u3�^]� �E�H�� UQj j �@0j j �u���   �uRjV�Ѓ�(^]� �����������U��Q�I��u3���]� � U�U�Rj j �@0j
jd�u�E�    ���   j �ujQ�ЋE���(��]� ���U��Q�I��u3���]� � U�U�Rj j �@0j
jdj8j �u�E�    ���   j	Q�ЋE���(��]� ����U��Q�I��u3���]� � U�U�Rj j �@0j
j j8j h�  �E�    ���   jQ�ЋE���(��]� ��U��Q�I��u3���]� � U�U�Rj j �@0j
j j�u�E�    �u���   jQ�ЋE���(��]� ���U��Q�I��u3���]� � U�U�Rj j �@0jj j?�u�E�    ���   h�  jQ�ЋE���(��]� �U��Q�I��u3���]� � U�U�Rj j �@0j
j �u�E�    �u���   �ujQ�ЋE���(��]� ��U��QV�q��u	3�^��]� �E�E�    �H�� UQ�M�Q�@0RV�@8�Ћ�����tK�U���tD� U�uR�A�@�ЋM�����t(� UQ�@�@�ЋM�����t� UQ�@� �Ѓ���^��]� �����������U��V�q��u3�^]� �E�H�� UQ�u�@0RV�@0�Ѓ�^]� �����������U��V�q��u3�^]� �E�H�� UQ�u�@0RV�@,�Ѓ�^]� �����������U��V�q��u3�^]� �E�H�� UQ�MQ�@0RV�@,�ЋM3҃�9U�^]� �������������U�� U��$�@Vj ��M܋@hCITb�С U�M��uhCITb�@�@8�С U�M�j hsirt�@�@4�С U�M�j hulav�@�@4�ЍE܋�P�u�E�P�H���� UP���   �@8�Ћ U�����E����   P�	�ы U���A�M܋@�Ћ�^��]� U�� U��$�@Vj ��M܋@htlfv�С U�M��E���@�$hulav�@,�С U�M�haerfhtmrf�@�@4�С U�M��E ���@�$hinim�@,�С U�M��E(���@�$hixam�@,�С U�M��E0���@�$hpets�@,�С U�M�j hsirt�@�@4���U8W�f.џ��Dz�E@f.����D{?� U�M܃��@�$h2nim�@,�С U�M��E@���@�$h2xam�@,�С U�M�j hdauq�@�@4�ЍE܋�P�u�E�P����� UP���   �@8�Ћ U�����E����   P�	�ы U���A�M܋@�Ћ�^��]�@ ������U�� U��$�@Vj ��M܋@htniv�С U�M��uhulav�@�@4�С U�M�hgnlfhtmrf�@�@4�С U�M��uhinim�@�@4�С U�M��uhixam�@�@4�С U�M��uhpets�@�@4�С U�M�j hsirt�@�@4�ЍE܋�P�u�E�P����� UP���   �@8�Ћ U�����E����   P�	�ы U���A�M܋@�Ћ�^��]�  �����U��Q��j jj �u�u�����Y]� ���U��V�q��u3�^]� �E�H�� UQ�u�@0RV�@�Ѓ�^]� �����������U��I��t'� Uj j j �@0j j j �u���   j jQ�Ѓ�(]� ����������̋I��u3�á UQ�@0�@�Ѓ�����̸   ����������̡ Uj j j �@0j j j ���   j j j4�q�Ѓ�(��������V��N��u3�^� � Uj j j �@0j j j ���   j h� jQ�С Uh�  h�  j��@0j�j j�v���   �Ѓ�D^� ��������������U�� UVW�}��@�ϋ@ ��=NIVb��   ��   =TCAbktA=$'  t'=MicM��   QhIicM���������WP�R_^]� ���W�P_�   ^]� � U��j hdiem�@���   �Ћ��WP�R_^]� =INIb��   �~ u�����F   �P_^]� �~ t�����P_^]� =atniHt1=ckhct=ytsdu?����P_�F    3�^]� ����P_^]� � U�@�@`��_3�^]� =cnyst_3�^]� � U��j hIicM�@���   �Ћ��WP�R_^]� ����������������������� �������������3��������������̸   � ��������V��N��9��t� UQ�@0�@�Ѓ��F    ^������̡ UV��Vh�� ��9�@0� �Ѓ��F�F    ��^����̡ Uj0Q�@�@@�Ѓ��������������U��(U��V���u[� UjhD �@���   �ЋЃ���tK� U�A�M�Q�M�Q���   �M�QR�Ѓ���t&�E���t�(U�xh|��t�@h��t	�uV�Ѓ�^��]� ������������U��(U��V���u[� UjhD �@���   �ЋЃ���tK� U�A�M�Q�M�Q���   �M�QR�Ѓ���t&�E���t�(U�xd|��t�@d��t	�uV�Ѓ�^��]� �����������̋ѹD h(U�  ��������������U��(U��V���u[� UjhD �@���   �ЋЃ���t\� U�A�M�Q�M�Q���   �M�QR�Ѓ���t7�E���t0�(U�x\|%��t!�@\��tV�Ѓ����u������u���2�����^��]� ���������U��(U��V���u[� UjhD �@���   �ЋЃ���tK� U�A�M�Q�M�Q���   �M�QR�Ѓ���t&�E���t�(U�xx|��t�@x��t	V�u�Ѓ���^��]� ����������U��(U��V���u[� UjhD �@���   �ЋЃ���tH� U�A�M�Q�M�Q���   �M�QR�Ѓ���t#�E���t�(U�x\|��t�@\��tV�Ѓ���^��]����������������U��(U��V���u[� UjhD �@���   �ЋЃ���tR� U�A�M�Q�M�Q���   �M�QR�Ѓ���t-�E���t&�(U�x\|��t�@\��tV�Ѓ����u������^��]� ���U��(U��V���u[� UjhD �@���   �ЋЃ���tH� U�A�M�Q�M�Q���   �M�QR�Ѓ���t#�E���t�(U�x`|��t�@`��tV�Ѓ�^��]��U��(U��V���u[� UjhD �@���   �ЋЃ���tg� U�A�M�Q�M�Q���   �M�QR�Ѓ���tB�E���t;�(U�x\|0��t,�@\��t%V�ЋE���E�΍E��E�    �E�    P�������^��]� ��������������U�� U���@Vj �u��X  ��M�hicMCQ�Ћ U���    �F    j ���   RV�@�С U�M�Q���   � �Ѓ� ��^��]��������̡ U�@��p  ��U���� U�U�R�U�R�@�U�RQ���   �Ѓ����#E���]���������������̡ UjQ�@���   �Ѓ����������̡ Uj�@�@,��Y���������������̡ U�@�@`����̡ URQ�@�@@�Ѓ���������������U�� Uh�   �u�u�@h� jh�>  ���   �Ѓ�]�̡ UQ�@�@��Y�U�� U��4�@V��p  �Ѕ���   � U�M�j h���@�@�С U�M�Vh���@�@4�С U�M�j h���@�@4�С U�M�j Q�M��@hicMCQ��X  �Ћ U���E�    �E�    j ���   �M�RQ�@�С U�M������   Q� �С U�M������   Q� �С U�M̃��@�@��^��]á Uj �@��D  ��Y�������������U�� U���@VW���M䋀�  jQ�Ћ U��W�I�I�ы UW�A$�@D�С UWV�@$�@L�С U�M�Q�@$�@H�С U�M�Q�@�@�Ѓ� ��_^��]����̡ UQ�@�@�Ѓ����������������U�� U���@$VWQ�@$�M�Q�Ћ U���}W�I�I�ы UW�A$�@D�С UWV�@$�@L�С U�H$�E�P�IH�ы U�E�P�I�I�у� ��_^��]� ���̡ UQ�@$�@�Ѓ����������������U�� U���@$VWQ�@�M�Q�Ћ U���}W�I�I�ы UWV�I�I�ы U�E�P�I�I�у���_^��]� ���U�� U�uQ�@$�@<�Ѓ�]� ����̡ UQ�@$�@h��Y�U���4�E�VWP����� UP�E�P�I$�A�Ћ U���}W�I�I�ы U���AWV�@�С U�M�Q�@�@�С U���H$�E�P�IH�ы U�EЃ��IP�I�у���_^��]� ��������������U�� U���@$VWQ�@ �M�Q�Ћ U���}W�I�I�ы UW�A$�@D�С UWV�@$�@L�С U�H$�E�P�IH�ы U�E�P�I�I�у� ��_^��]� ����U�� UV��V�@�@�С UV�@$�@D�С U�uV�@$�@�Ѓ���^]� ���U���<SV���E�    �8UW��t�EĻ   P�������-� U�M�Q�   �@�@�С U�M�Q�@$�@D�Ѓ��}� UV�@�@�С UV�@$�@D�С UVW�@$�@L�Ѓ���t(� U�M�Q����@$�@H�С U�M�Q�@�@�Ѓ���t%� U�M�Q�@$�@H�С U�M�Q�@�@�Ѓ�_��^[��]��������U�� U���@VW���M�@$Q�Ћ U��W�I�I�ы UW�A$�@D�С UWV�@$�@L�С U�M�Q�@$�@H�С U�M�Q�@�@�Ѓ���_^��]���������̡ U�@�@�����U�� U�@�E   �E� � ]���̡ UV��V�@���   �Ѓ��    ^�̡ U�@���   ��U�� U�@���   ]��������������U�� U�@���   ]��������������U�� U�@�@|]�����������������U�� U�@�@p]�����������������U�� U�@�@L]�����������������U�� U�@�@,]����������������̡ UQ�$�@�@$���������������U�� U�@�@]����������������̡ URQ�@�@�Ѓ���������������U�� UV��V�@$�u�@L�Ѓ���^]� ��������������̡ UV��V�@�@�С UV�@$�@D�Ѓ���^�����������U�� UV��V�@�@�С UV�@$�@D�С U�uV�@$�@d�Ѓ���^]� ���U�� UVW����@W�@�С UW�@$�@D�С UWV�@$�@L�С U�uW�@$�@@�Ѓ���_^]���V���������^�����U����E�VP���>���� U�M�Q�@$�@�Ѓ���tY� U�M�jQ�@�@�Ѓ���u�M�������t3� UjV�@�@�Ѓ���u� UV�@�@�Ѓ���t�   �3�� U�H$�E�P�IH�ы U�E�P�I�I�у���^��]��������������̡ UV��V�@$�@H�С UV�@�@�Ѓ�^�������������U�� UV��V�@�@�С UV�@$�@D�С UV�u�@$�@L�Ѓ���^]� ���U�� U�uR�@Q���  �Ѓ�]����U�� U�u�u�@RQ��  �Ѓ�]�V����t� UQ�@� �Ѓ��    ^����������������U�� U�uR�@Q���   �Ѓ�]����V����t� UQ�@@�@�Ѓ��    ^��������������̡ Uh���@@���   �Ѓ���������U�� U���   �E    �@ ]�������U�� U���   �E    �@]�������U�� UV�u��@j��@�Ћ�^]� �U�� UVj �u�@��@�Ћ�^]� �U�� UVj ��M�@j V���   �Ћ�^]� ����������̡ U�@�@����̡ UVj j��@��@�Ћ�^���������h,U��   �/D �  �����������U��,U��V���u^� Ujh/D �@���   �ЋЃ���tX� U�A�M�Q�M�Q���   �M�QR�Ѓ���t3�E���t,�,U�x�   |��t���   ��t�u��j ��^��]� 3�^��]� �������������U�� UV��@l�v�@�ЋM����u�A^]� � U�u�u�@lQ�u� ��3ɉF��������^]� �������������̡ U�q�H:�@l�@��Y��������̡ UV��@@�6�@�Ѓ��    ^���̡ UQ�@H� �Ѓ�����������������U��E��HV���2  �$���   ^��]á�U@��U���  �E� U�8�>  }
�����^��]Ëu��t�U��E�P:�   �E�M   �E�    �t�������   ���5����Љ8U����   � URV�A$�@L�Ѓ��   ^��]ËM������^���H��]�������^��؋�]���UuW�F  ������58U��tC� UV�@$�@H�С UV�@�@�Ћ8U����t� UQ�@� �Ѓ��8U    �   ^��]Ã��^��]Ë�e[����������U���Mu�E�4U�E�0U�   ]� ��������������̃y ��:u� U�q�@P�@��Y���U��M�]�`����U��M�]�`����U��M�]�`���̋I��t� UjQ�@P�@�Ѓ�� ���� ���������U���V�uW����t���u]� UjQ�@���   �Ћȃ���t?� U�UR�U�R�@�U�RQ���   �Ѓ���t�E��t��t�3�;x_O�^��]�3�_^��]�������V����t� UQ�@� �Ѓ��    ^����������������U��M�US�]V3�W�}95�U~(�d$ ��UWSQ��R�Ѓ���u!�MF�U;5�U|�WSQR�DU��_^[]�_^�   []Ë�U��t� UQ�@� �Ѓ���U    ��U    ��U    ���%x Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ����%| �%� �������̸@A������������������������̋�U��t� UQ�@� �Ѓ���U    ��U    ��U    �                                                                                                                                                                                       nD XD BD (D D D �C �D     �B �B �B �B C C "C *C �B BC PC ZC nC �C �C �C �C �B �B 4C �B �D �D �D                      " �!             ���Y       �   (; (/     ���Y          �; �/ �;�      RPR    }Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������-DT�!	@}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������       }Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I��}Ô%�I�T}Ô%�I�����������������}Ô%�I�T���������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I��       �����������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������}Ô%�I�T}Ô%�I���������}Ô%�I�T}Ô%�I�������������������������$filepath$filename_$pass    No object ID found   Object(s) ID Added Done,       c:\program files\maxon\cinema 4d r16\plugins\easyobjectid\source\maincommand.cpp    Easy Object ID v2   �<� �� � �� ` �� �� �  � �� p� @< � �  � �   �� �� �� � �� p� ?� �� � �� 0 �� �� � @� �� p� >�  � � Ь � �� � � �� �� p� �>� �� � �� � �� �� � �� �� p� �=� � � � � �� � � � �� p� �=�� � @� � � �� �� P~ � �� p� D>0 �(  � p( `( �� �� �� �� p<� �c �^ ��\ ���PEasyObjectId    plugins Configuration.data  EasyObject ID v2 - Settings     Vray Settings   Consider For AA Affect Matte Object Octane Settings Define Object ID    Define Layer ID Redshift Settings   Reflect/Refract IDs Multi-Pass Output   Enable  Bits Pers Channels  8 Bits  16 Bits 32 Bits File Output Path    Data Type   RGB RGBA    Format  OpenEXR TIFF    PNG TARGA   JPEG    Half Float (16 Bits)    Float (32 Bits) Compression None    Default LZW CCITT RLE   ZIP PackBits    RLE ZIPS    PIZ PXR24   B44 DWAA    DWBB    DWA Compression JPEG Compression    Storage Scanline    Tiled   Ok  c:\program files\maxon\cinema 4d r16\frameworks\cinema.framework\source\c4d_misc\datastructures\basearray.h Object Buffer Driver    ObjectBuffer_       E'  '.*L    Oject_ID_   modules resource    res c:\program files\maxon\cinema 4d r16\frameworks\cinema.framework\source\c4d_resource.cpp    T?0 �?� ��� ��� ���Ph?� �� p� �� ��  �  � �� �� �� �� �?@ �c:\program files\maxon\cinema 4d r16\frameworks\cinema.framework\source\c4d_pmain.cpp   @� � � �      �Ngm���         �Ngm��C      �?H                                                           P        RSDS��]ӗ@kJ����C��   C:\Program Files\MAXON\CINEMA 4D R16\plugins\EasyObjectID\_obj\EasyObjectID\Win32_Release\EasyObjectID.pdb      5                          P�;           �;�;    P        ����    @   �;           >�==    dP       ����    @   p=            �P�>�P       ����    @   =            �P�>�P       ����    @   �=            �P=�P       ����    @   �=�P       ����    @   �>�<(>    L==               H?@P        ����    @   �=0Q       ����    @   ?�P       ����    @   �>=               X>           �>            @P�=�<t>    pQ       ����    @   d>            �P�=           h=,?=               �=t>                LQ�>Q        ����    @   �>            0Q?$<=               <(P        ����    @   <           �<�<=    (>               �>            dPp=           �<0=�<t>               �=            pQd>           �>LQ       ����    @   �>T<=                (P<            �Q�?�?               |?            Q�>�Q        ����    @   �?�?               �?�Q        ����    @   �?            �Q�?            �QD@�Q        ����    @   D@ @               <@                    ����    ����    ����    �!     x! �! ����    ����    ����    �"     ����    ����    ����    #     ����    ����    ����G# p#     ����    ����    ����y$ �$     �Qx���o� ����    ����                  A"�   A   ,A                                ���Y    �A          �A �A �A @ �A   EasyObjectID.cdl c4d_main B         �B $  �A         �D                        nD XD BD (D D D �C �D     �B �B �B �B C C "C *C �B BC PC ZC nC �C �C �C �C �B �B 4C �B �D �D �D     I_purecall r ??3@YAXPAX@Z  p ??2@YAPAXI@Z  �free  MSVCR120.dll  o ??1type_info@@UAE@XZ  o__CppXcptFilter _amsg_exit  �_malloc_crt _initterm _initterm_e �_lock _unlock ._calloc_crt �__dllonexit :_onexit 5?terminate@@YAXXZ �__clean_type_info_names_internal  z_except_handler4_common P_crt_debugger_hook  �__crtUnhandledException �__crtTerminateProcess gIsDebuggerPresent !EncodePointer � DecodePointer -QueryPerformanceCounter 
GetCurrentProcessId GetCurrentThreadId  �GetSystemTimeAsFileTime mIsProcessorFeaturePresent KERNEL32.dll  t__CxxFrameHandler3  �memcpy  �memset                                                                                                                                                                                                                                                                                                      ����N�@���D    �     .?AVtype_info@@ �     .?AVBaseData@@  �     .?AVDefaultRenderManager@@  �     .?AVVrayRenderEngine@@  �     .?AVArnoldRenderEngine@@    �     .?AVUi@@    �     .?AVCommandData@@   �     .?AVC4DRenderEngine@@   �     .?AVIrayRenderEngine@@  �     .?AVGeDialog@@  �     .?AVMainCommand@@   �     .?AVOctaneRenderEngine@@    �     .?AVRedshiftRenderEngine@@  �     .H  �     .?AVGeUserArea@@    �     .?AVNeighbor@@  �     .?AVC4DThread@@                                         �                  0  �               	  H   `` }                  <?xml version='1.0' encoding='UTF-8' standalone='yes'?>
<assembly xmlns='urn:schemas-microsoft-com:asm.v1' manifestVersion='1.0'>
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level='asInvoker' uiAccess='false' />
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>
                                        000!010d0u0�0�0�0n1w122d2n2t2�23$373E3W3h3v3�3�3�344434<4h4t4�4�4�4�4�455#5R5�5�5�5�5"6�6�6�6�6�647=7X7�7�7�7D8v8�8�89q9v9:!:^:�:�:�:);7;I;~;�;�;�;<<E<�<�<�<�<�<=+=D=P=h=�=�=�=�=�=�=*>4>9>>>T>`>�>�>�>�>�>�>�>�>??'?1?7???o?w?|?�?�?�?�?�?�?�?�?      X  00!00080O0U0�0�0�0�011c1�1�1�1�1�1�1�1	22"272B2X2r2|2�2'3�3�3�3�3�34+4?4E4�455&5/5<5k5s5�5�5�5�5�5�5�5�5�5I6N6^6d6j6p6v6|6�6�6�6�6�6�6�6�6�67777!7(7/767>7F7N7Z7c7h7n7x7�7�7�7�7�7�7�7�7�788�8'9l9}9�9�9�9�9�9::):@:U:f:z:�:�:�:�:�:�:�:;*;C;V;g;{;�;�;�;,<=<O<Z<m<�<�<�<�<�< ==&=:=L=W=h=�=�=�=�=�=�=>>'>;>O>c>�>�>�>T?�?�?   0  8  0_0�0�0�001~1�1�12"272\2�2�2�2�2�2�2�23#3G3U3g3z3�3�3�3�3�3474Z4r4�4�4�4�4�45/5J5e5�5�5�5�5�5�5606J6\6�6�6�6�67)7G7e7x7�7
8D8^8o8w8�8�8�8�8�8�8�899(999Q9f9x9�9�9�9�9�9�9�9::(:?:S:^:l:�:�:�:�:�:�:�:�:;;*;B;S;d;y;�;�;�;�;�;�;	<<+<<<M<^<r<�<�<�<�<�<�<=0=_=|=�=�=�=>->U>}>�>�>�>?E?m?�?�?�?   @  �   050]0�0�0�0�01)1i1�1�1�1�122@2Z2�2�2�2�24;4`4�4�4�4�45.5Y5�5�5�56L6t6�6�6 7(7d7�7�7�7858]8�8�8�89+9`9d9h9l9p9�9�9�9:A:U:j::�:�:�:�:;0;�;�;�;�;�;#<4<K<`<u<�<�<�<�<�<=n=�=�=�=�=>>.>C>X>�>�>�>�>�>	??4?I?^?�?�?�?�?�? P  �   00.0C0X0�0�011*1?1j1{1�1�1�1�122[2l2~2�2�2�2�2�23>3R3i3~3�3�3�3�344J4^4u4�4�4�4�4�45%5V5j5�5�5�5�5�56616b6v6�6�6�6�6�67(7=7�7�7848e8�8�8�8)9U9�9�9:9:e:�:�:�:;P;|;�;�;<8<i<�<�<�=>>>>>   `  �   �2�2�3 44%4N4`4r44�4�4�45$515M5�5�5�5�5�5�566;6W6h6z6�6�6�6�67797K7]7j7�7�7�7�7�7�7,8I8[8h8�8�8�8�8�8�8�89.9I9[9h9�9�9�9�9�9#:K:u:�:�:�:�: ;$;A;k;�;�;�;�;<9<K<|<�<�<�<�<=%===O=\=j=�=�=�=�=�=	>(>R>|>�>�>�>�>?1?U?r?�?�?�?�? p  �   050_00�0�0�0�0-1?1p1�1�1�1�1202T2�2�2�2�233N3`3�3�3�3�34.4Q4u4�4�4�4�4,5>5o5�5�5�5�56=6O6r6�6�6�6
77M7_7�7�7�7�78(8\8n8�8�8�8�8.9@9t9�9�9�9 ::F:c:�:�:�:�:;/;Y;y;�;�;�;�;%<E<i<{<�<�<�<=6=`=x=�=�=�=�=�=>/>�>�>�>�>?N?n?�?�?�?�?   �  �   00J0�0�0�0�0 1 1=1a1o1�1�1�12?2M2_2�2�2�2�23$353A3O3h3�3�3�3�3Q4�4�4�4�4�45U5o5x5�5�5�56%6@6Y6n6�6�6�6�6�6�677,7A7Y7�7�78*838T8�8�8�8�8�89F9f9�9�9�9^<x<�<�<�<�<=<=v=�=�=�=>(>c>�>x?�?�? �  �   090J0e00�0�0�0181Q1�1"2M2k2�23-3Q3z3�3�3�34<4Z4�4�4�455(5I5x5�5�5�5�5;6_6�6�6727;7\7�7�7�7�78-8Z8c8�8�8�8�8�8)9H9�9�9�9�9�9�9:;:c:}:�:�:�:�:;.;�;�;�;�; <<:<V<�<�<�<�<=)=9=O=g=|=�=�=�=�=�=>->O>l>�>�>�>�>�>�> ? ?4?H?]?p?�?�? �  �   �0�0�0�01.1B1Z1p1{1�1�1�1�1�1�12282M2k2�2�2�2�2 33$3E3w3�3�3�34r4�4�4�4�45E5e5�5�5�5�56!6F6T6m6�6�6�6�667Y77�7�7�78'8X8a8�8�8�89,9[9�9�9�9�9�9:8:O:�:�:�:�:;;4;F;�;<*<6<W<�<�<=4===^=�=�=�=�=U>x>�>�>?1?e?�?�?�? �  �   0>0G0l0�0�0�01A1f1�1�1�1�1�1252n2�2�2�2 3+3>3J3k3�3�3�344�4�425|5�5�5�5�5636]6�6�6�6:7\7e7�7�7�7�7;8\8�8�8�8�89W9w9�9::@:u:�:;0;9;Z;�;�;,<J<S<t<�<�<�<=)=B=W=�=�=�=>R>t>}>�>�>�>?�?�?�?�?   �  �   0�0�0�0�0�0)1�1�1�1�12<2�2�2�2�2-3P3t3�3�3474@4a4�4�4�4K5i5r5�5�5�5_6}6�6�6�67y7�7�7�7�78�8�8�8�8939�9�9�9�9+:N:�:�:�:
;?;b;�;�; <!<V<y<�<�<+=T=�=�=�>�>�>�>$?G?�?�?   �  �   /0�0�0101T1p1�1�1�1�12!252L2c2z2�2�23C3f3�3�3�3#474h4q4�4�4�45<5k5�5�5�5�56'6H6_6�6�6�67+7B7a7v7�7�7!8;8S8x8�8�8�8�8�8�8	9#989V9m99�9�9�9::8:j:�:�:�:�:;J;�;�;�;�;�;'<f<�<�<�<�<=/=f=}=�=�=�=�=>>5>M>}>�>�>?&?G?v?�?�?�?�? �  <  0>0^0z0�0�0�0!1D1i1�1�1�1(212V2�2�2�2�2+3P3n3w3�3�3�344X4{4�4�4�4555Q5Z5{5�5�5�5�56>6S6{6�6�6�6�6
717F7d7v7�7�7�7�7�7�78 818<8H8Z8f8�8�8�89"979T9f9�9�9�9�9�9::,:B:T:i:x:�:�:�:�:�:�:�:;(;=;U;r;�;�;�;�;�;�;<<.<F<^<s<�<�<�<�<�<�<=4=C=[=l=}=�=�=�=�=�=>>$>*><>G>P>^>m>y>�>�>�>�>�>�>�>?4?N?b?r?�?   �  �   0!0D0q0�0�0|1�1�1�1�1�1�1�1�1�122%2�2�2�3�3�34�4�4�4-5a5{5�5�56#6�6$7?7�7�7�78)808d8�8	9�9�9�9�9J:h:�:�:�:�:A;S;k;�;�;�;�;<=<<�<�<=M=�=�=$>t>�>?d?�?     �   0:0U0m0�0�0+1d1�1�1�1�1�12$2A2c2}2�2�2�2383Z3�3�3�3�3�3	4#4;4S4k4�4�4�45K5�5�5�56T6�6_7�7�78!8*808Q8t8�8�8�89949_9�9�9�9�9:T:c:�:�:�:�:;?;t;�;�;�;<<4<_<�<�<�<�<4=Y=|=�=�=�=>1>A>d>�>�>�>�>�>?&?M?c?y?�?�?�?�?�?    8   0010T0l0�0�0�0�0�0�01 101T1q1�1�1�1�1�1�1$2<2P2^2m22�2�2�2�23%3<3J3X3o3�3�3�3�3�3�344,4Q4d4�4�4�4�4�4545T5q5�5�5�56646E6S6t6�6�6�6�6�6!787V7h7�7�7�7�7�78$8J8t8�8�8�89$9D9d9�9�9�9�9�9:?:�:�:�:�:;!;W;f;l;};�;�;�;<1<:<H<W<c<t<�<�<�<�<�<�<�<�<�<�<8=R=x=�=�=&>1>N>Z>r>{>�>�>�>�>�>�>�>??,?6?@?      �0�0�0�0�0�0�0�0�0   0 �  �4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:�:�:�:�:�:;�;�;�;�;�;<<<<$<<<L<P<T<l<|<�<�<�<�<�<�<�<�<�<�<�<�<�<==,=0=H=L=d=h=|=�=�=�=�=�=�=�=�=�=�=�=�=>> >$>(>@>P>T>X>\>p>t>�>�>�>�>�>�>�>�>�>�>�>�>???(?,?D?H?L?`?d?t?x?|?�?�?�?�?�?�?�?�?�?   @ 4   0000 080<0P0�0�0�0�0�0�0�01111<1H1P1 P ,   0(0@0d0�0�0�0�0�0101L1p1�1�1�1�1                                                                                                                                                                                                                                                                                                                                      